BZh91AY&SY���� ߀Py���g߰����`
=�����  A� $����@P    5=�����bmG�`A�hbi�4d1?O�S@�@    M$�Ҧ��1D� h sFLL LFi�#ɀFI &�0�i�m'����Sa=M�='Ꞧ�Г�u�$Db�3~u9)tD�	K�ϝ��%��,T%�"T�q'�Jә�	' n��B@WЕ,TJNUrR4��� � ZS31̹�q��2�s2�c[h����n9���e�g��73���)���w���ޑ`��ۻN��<�-Ӧx�x÷F�����Ӣ	��P��dL��=��c-E	dqC��.��3�g���=?��=�C��C|�C�I*��o���H-^J��D��g��yqV�I�3�zG脄�V�1x�v�Ln�0����I�3�X:����/.���I/.�E����P4j��[ ,�k��@$�+{<��#9���ff'�ɡ�Z�p�A@�	_�J@������{�ns��?�Q��]�Sb��DKr�C=�d�=�6���k�%��:c"[���uN5
�!�CC��m�]���0�gV�>#�a�H�E�a�u4�E�>�o��
�M��	�l!S	<l�c�ia�iφ�{Z�m�z���C������(�0�Hp+���� ,����٤E9P��~�?HdxH�4n�Y �r��T�4�>���Y�,t��D@s�M��3�"�50Z�Q0�Q
��Q���@�ف���[�����|{����}�s�Ӱ�ݺ���*J�Q4o�/.�ۑx�&�z3^F�f���*r��,<pp0х��w�ζ�����&$�b6�~�C�D�8yS0l'Tx�OL�q��4�(�;�xԲk%ėe��׸gR�����1]�OgC�Y$����;�����yWX�/֡-[�1��S�䑆9�|7͠ClP��2�hC�L�ԗH{�0I$�y'1�f�Y0�-���-z(�����m�|R0E��F^rS���80ipC'i��TI$ξf�Q4�uyn���j�5�+mw��-�4�� C兠B`;�є����by������롶�	������ɰ�0�3��\�f��Sf�P;���X*��	T�Ӷ*L�CMG&�3�`��0˻�j`�Ϙ��=4�����~��#��t׃�X���,DD_

�d������N�N_��\��O�E(�Ȑ16��#D ��h2 �A�K`Y$�Y79�Ѥ��G00�Id���%Ė�d�iNѹd�3fi��R�AT��<�mo+��g��<�iv0x[q{���p8�iw�X �%��3g��97�i��mr�Ӭ��Z�7b��{S�|R��o{�ѣ�L[]1"v&o����_���9���RH�ܴ)E��L�Oj���8��O���n�y�>��OT��џ�H��&=&כ�>=�Nѣ����Qd�'d֎D�xJY��NX,*�v��V�pN�Iz���\޾���^8j�p�>�/	ܨ�4��WW	�=���R�g�}�6Gw�jL&��-ER"�(T�*�Yf��2�[�u�|!T�ӹ��M��KҖLKc�"��)�Z�3�c�,TH�83Z�n�f?ze�=,%<�`�+<8N�׬�8�O�0+�(��Of\ZӔH�4p�+�^��{a�qN4I'�;�0�º��ϩuNl#7b��N%���_;c����{��%��m�k������~��b�5�_�ד�ZA�0�Sܢڔ�kTb|		-%�;.�.J�qr�ĸ�������|waű,M�l����[g'S9N����%���_7k'0Ԓ8�;�l��pUQEUQEUTQTUQUUUUUQQUUUUTTQUPUUE}�x6� S+��md�Gc�{P�T̖��ժ]�tT�s�u�,�9i��L:�3�c%��L'S���bD����ѻ)X��r3�̜�K&�N2��ɛ90w*�0%�{�a�9����}�؇�혷�p�b���d��
�G~_.��b��g�'�rE8P�����