BZh91AY&SY'ޠH �_�@y���g߰����`��K � �8��TRPI"i�	�B�M���ښdhh�44�hE=��JQ	�	��F�	��@������10 &M4hѦA�0�!��&@�M     i��&�&	��0`��"HD���S�1Oj���=@0�M���(Ay�@���D�p����	���|�.Q�(�tQ��A��(�.�1\��|
�eSw?F�=���� &	I � 	 " � ! �$�|��uT�!{�YZ�(@yy�6]�_%jdDhLдh��4$�(�ta�,�e;�1�/��"�de��5f/�-���4��')���y]c�&�3��<��!�J�቞!  ���<�'um�m=�V5���K$�D$�+I�bH��DE$�����%I%�H2I$��IDD$��L���		���m[G�<:��3�,xo�CK�q��H�uy�`2�c�$��z�h�i�<��������Z��Z]M!2����T@�N0�m��@Uj��Z�a�6���j�F1��L��T�Fn A	B&�%�)�+Zc8���o8gp��H:v1��+l�a.��m�w"t�&Xh�Gr#
PZ6����P��,���!t �����lH7��q��F��m��[��1Ӧ�����Ƶ��Nr_ YoGJץR������YkQ|+�%��m�[2�5�&s�Ί�|7����.�j�^��S�$���.b��9!��   ��M����^I��ȔԗFQc�6�v;(��=�<D;9���    =�)�k���������Ⱥ6F�y�vs���k�p  K̴�|��ݦӲd�h��k�fU5����C��J���'�u����y����&����X�7*���S�a �Ϛq��6����)��F����{��Lз�����E�Y�q4X8��wz8�c���㤑��$��$�4Q���{�3�т�c��]w��l��0!�h#0 x���#U ��"@�$� ���j]*�iok�T
((�(&p�ST1�KM^���{{JI@�_��o�c�J"Q���:3t��U�K���Η�ώ��]\JxI�&���b�gq}�s��0�GY��)1��Є�ģ�7[�A�]���-
?���z����!9�=�,�E��x�4�w�iԄ�1����."\�\*K��a��)�e���
(�5hr⑱('I�Lm/9(4�qx�N��; ������ #jڴ�~��F�Qc��c̞[��)�$`���|��`��u�Y,�P^�&"(�-9S��k��|��ȣc��ʥ��}'N^�?#���<�̰�tgZQ+:��&f���m�=A�Ʃd����<a�m�+�w��_�;Y�LL�V��9x�`����ټo�V]�}�[!G����PBk*Oi���a�ƨn#Z�hZ�>F���4����o7����o��ia�8S����!��b��[��tt8���78�:(J=G[wf��\̈�F�u1�1��r����42�YÚt�t��js�8Sҋ�C&�`=ٜhW�G}���qD�m���A���kԧBB����0��0'��H���Ƈ�32��C���>eě�V�a1*Pw1�L]#"8b��3+���H�!��;�+��]��B@�z� 