BZh91AY&SY
 �_�@yc���g߰����`�\�yU��P ��jCɑ�hA�4M�@5= �U<��� A�4h  jm�IOԀz�i�� ��  $$@�Pd ��dh    ���a2dɑ��4�# C T�j4��&L����M@i��	;!R�S�x����$�D���ؖ��z�"%L�=����U����$Т1�OE%�LhΞ]~N���     �   A �� @ m�p�{����0���6�۱{eE�R��&�[]뒥Vb���R�sjޚ"&��1�C�2�$(��:� �F˫�
X�]8|oh��gŭ�5(�M�G3	E�$����=Z�%7�ͫ.�s]�O8��*cq"㎒8�@D�|X&B>��i��-J��4�M�ISHݬ̰��Jg*�2�k��I*���ř���:I:J���{��;��*
"�V���B��Ud;-�:��
]Ul���� ��`��!�b�$ͫD֑eJۺzF��C\���`��f�4gzd�i_�Mhi�!���;iWJ���а��MZՁ�5�ƢFrb��i2���@��E�a Q�N�$�8@y�r	�fN��_C��ߖ��Ǖ��a���j���Ս���'\ӫ8r뇏,�s��c^oq�uZ�o'�Y�����i���RZ`͒�݂�m ��A���l�PMfMU�qN�rv�"�8��.�S;=o�D!R�Q�A��:� �H��؋�]��0�*�de��(S�%l�%Z5���kR�^�	��O.�]��O23�S@ͽ��� f�8�0�;a�uCd H$#_�C4�f��u�K͋S����
j�}���� �LJ�12w���K�#����ky�do� �c�Q�g�P���@�I��v՞n�w���cTI�������m�d��I��9">�ZH�*���w���m�)u[�;C��;c� x��@c�|M���!B.< ��bvU)~;�7X�'DSň�ƨ
N1B���40i0hi�S 4�/)\p�EL
("bĠ��SR����(K&U�T34ՋQ&kC��M ��M���g��$��s>L��?I��^����>V*�q�@0�I�~�AӚ�i�� T�O���^D�(���Br�s�f3G詋��H��f��W�����F���~�4�R"E�a�k>5>w7 ���9R����,��?�<Q����D�IŖ����wz0��#'��$�(�؇�6����z:pZ�Y+��Z��rx2/V�M��Z2�ޜ3z���_!�P��Qu�� 5���"��gP��?\+1X4�D��RAR�Jm켎��Lg��i摮j�U7�B�|�ǁ�y���)-t�]ˇl��vy��f���S�b�+�*|���D�p0�iz`��5{�v�'D��7U%c�a~Âj7�hI:���
�u:���z�:0�5s�7����a��0�JL'����I(�k@a���
�A��Y2(߹;��(��5O�3��I�zS ���U��_/>શ��<���5��e����f��p�冾ދ�.5T�Y�ȧ��<VIg�<e�C�g/��isI�u:^i�3����/3jF��9k-m��,V��u��q6���k�w&Z'Nɞ<�%���~<܌Q)��kc�-j���-���Qhqb�İ��g3LX�����Z'��$���m�S�Md���&ɩ�h����X�t��F�	�_�~�ӽh�L%�6����"�(HwGW 