BZh91AY&SYW�bP �_�@y���g߰����`�5�AP* I5O�OI�Қ��h���bhhɠ��5O�JT�F�P24  � 2���&	�M0&!��& �F L�*j       i��&�&	��0`��"HD���ѓ)�#L�2hz��(|"�@K��9�a`�$���(�d(��(+u�� ��w�]�DC�zD2��������,X D�  �0��"2   �#�]B����1с���"�D�6D9�Y54<y�w�C)ݼY++�Ac�Y�Yn��1FS7a�b��`�vkb:���5_����ƔiH������ʓ0�yȽ��J�a�
V�Ռ ��_g^|vV{�|9��F��*e�ݶ����[n""�j��m�m�[s��m����s32�W^O$���00ͫ�N� �u������F�E9O��wu᱗��Ei$�U����I6q�!N��{Z��ְ�4�l��`lN��,'I$)B��0�dY��-��$C��ڲ�ɢ���!����M����#O`4
��R��:G������:T��[׌%�$RIw�~@FZI�[	0�{0��L8a+&sqd�X�&�l��T��{߀ҙX�x��lZ�nQֺ�ً��I!�g����C���(w�U�-F�����6g{��0mf'x���Q�I$�N1gU9�������d�g�j&`VU99=�j虉&;̝�R�I$�[�lL��bDF���|���e�a�k:.s�6�Ġa��I$��&^�����qn�<BDdLe=��3��Ý�����̺ظ;��Y���=kK`��c�x;��c��@�v�TT�!x7��M��<U�'�|��l��ؕ�U�ǜ�H���-UY��;�vΞN��NA$�$�(qd��7vkZ���97{��"F��H1e��y_EgsFU���]���l��03���$�1�W�"@��AT� @�H�h��.ՠ�g^�fTh��
�ABj��Ii�ނ�8����S"$�� ����*.����F��^~~��΢��9�*?.\���~���f轩���w��(9��>a����1,&11�B�������芬��_��P�=ol��k�'N���dX�Wć@v8�:�7�	��/8�'��I���2$ �O,�V����V�F)�u��&{M�٩Ľ��Z4����}س��S��pm\��F�Q������c�>Ɓ�%��0�epL�S$��+����5pdt7�f8+��v�����ٗ3AF���*��:��\�s8�0.e�8����9�C������O�חa�Dlr:�	������T^
#�y���WQ�.^�ۄ��G#yb��Q���pG�n�6V^;_?G�Q�06u�J*Oi��v���T;�ք7�O��=A���`	G_����J�6(����^@���q�~�arqt�˓mD�ި��7(��E���ݬu3"�Ѡ�c�s�N���)�C*%�9�YwN@0H���s6\����Z���w�s9��K�L�n�L��f��|�.J#��n6��!�˔���h|9���;2!!���>eħ�̤�b6 �c�R_n��1����̰T��'�`5&�Wt��H�

�LJ 