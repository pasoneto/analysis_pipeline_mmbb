BZh91AY&SY�`8b �߀@y���g߰����`�z�x���T '#�f ��P���)�z�4�2&� �h�S�LԐ�h�	��& M4�b��������4ɀ #!��$$A2SF�4�  d 9�&L�0�&&��!�0# T�4A1�	�M��4�Ѡ z�5a�I��II�~, ��	���f�Q�?c@�!	�Z? ^�UU�1M%��|��Q/F�yz�vr�z�5   �  FE )  
uR�{��vhx�G+�\��Yf4��tZ�@t���P�����7�U�,)���F8؜�S�;�2�TU�,�m��(��A��'���n*V����~�$�ކ�?�֣]��\�Z���T����z!��T�����^��Z�a#� G��3�K0���x����s33��-���6�DCd��m�ݶ�n"!��m��m���C[�G��444tL��k$_��1��b�d]�m7��_������H�� �Ϩ$�T8�#������%�zW����̫�R�T��<�.6��}����wUe���e��h��XԼyƆ�͚0r=I��r������}LT��ոGbJ���-::����K:�>O-hZk��-/�a�ٮ��$�H��P#Y4$wS(l��A�mhM�QУ� �S}@1z4d0���j0��cv�ɍ_**ڈ^/�8ߺ�k��I$A�}��p��Wwz]�^��E77*E.�Mrk�m>�CU�k��69U�M$�I`�'P���$�
���&"�`@a_68�e��073;�l�;�$�I$��V�*$���$���z��(��/�Y��7��[MȡWi$�JE]
����OfT�.����(�8*�^B�sG��[��R)s=D�r�}���J����g�����TDy�Ҡs+#"Q�ed�O/�b*�[]XIt/��cldsw@�V)�-�3�� Q$�.�D��m�N@���̉U�������K�g<�x���1�i�&�m�А���9"18BU)~9pX�'F*ĥ�gh�EQS¬TQR�(����XZ(�����*(�`���9�E��`��b�Ӫ
N1LFZ�

��HY2�C3MX�av�q7��lHCi&�h5|�M�}Mt���f䊁��m?�$V��H{ٴTϯȇW�jmp�a_:�ZT�i���0�&r�c���X��=%yQ�~�c��i��H�����c�k���%L"ZG�G���#MUc3�B�+�Y	�IlMe�I�}�ƔP7U��y�j(��Y�{�I�=�vg�l�|�.>�E���F\�w�{���CZ��2���-�E��-ub��۱��?[&��wMI��$���R�J(�jg�Iy�-�{dsMʣK��c
hſ��fܺ"�"'s��3Z���|�{����yN9�L��q���t�z���^}	�]9���[�jN��L�J�?���;�	�j8T$��􊑾���{
7^M
�d�a(m0;e��9Iy��I(��p|�[�b�Pd�f�7�N���h�|��F-�M֩2Ob\$�ĕgo����
�p�Q�`9M���������f�l�,i`6p�����Ud������T�K=󑉷X�1���B�<n/�x��r�.i�Y]�F��W5kFR��[�@��&'
ӛ[U�)��B	\(N,�>�Bоd���>n�$D�s����1�-S�e���J-��Xu�3���%S�sJ�O��&>��m
�5$�r1��8�2j����*:&9~�IR<��$ѯ7�.�p�!j�p�