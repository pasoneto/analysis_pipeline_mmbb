BZh91AY&SY��� P_�Py���g߰����`	?z���Y��  ]S�݀ �M'��M�d��    4 � I
iM0��0�20&O�U@ �� �d  	4�ҞB���њ�LF� M �A�101��&$@�h�������F���F������		?.�!hH��A�|�Ť$�B&=ߡ�`B��C(�Z*�3�8�&���T�{�,�eF�yws��:�o��iZ��m)ioF-���qq�A�" (
� � ��UgwUus��4o����gO�z�����Ǳ�t�(3���U�hU����DB��F�)�f��)X|��?b�\u`J=����B�e4���W�~]�������32;
���η�1�͛�-n�ӻ���:��k�)�U��e��M�4y�����+/��H�ñ�#��+�N���+���&��\Z������q\�%s�W��t˜i�+�ӯ���:�!$G�����@�iBF4�#
vr� @u*^��X����A8���#\-�u�`��%�E���Yx,�ad���W�w;��Tӷ[�]g��$�r�-��;\b��q]��1,�+��K{�7����`-FB���o8�o�)�I�G��q�x��!:�'L-�}?�����Q��)Y|�ks1֚l�1�r#��T`RD�"A�xJ��ذ����0 Շ���U-��J�=��\\�<
�<?a.:U~��Jy�R��ۦ5$2d���
�pL�5���X.p�Uc��^�����u�_��jl��˥Hb�*�2�j��W�fy�JFDV�y]-T��q�:��1`fc���7U�Kp#Bֿ*�.g�(cV��$�$ �'U���,@��H�8��l��1
�յ�bZ����|y�-0�mm)��K�i�3�j�6��s��I"��UD�~�n})��J�E�6R��"�uk��Q��'U�=�R�����^ �rd�0�d�c�L�&
Nؘ�W(�* �&�͜��	�/��]���'4E3��kx������PDF/ܪ���w�~��h��Y���~�՞--*엗�K�$:RJ�A0�mH6�\��k�E����Iz^��q0�Е�	Bl�D�3I���!�p�b$)"�U����+���m��ۛ�ÿ�N�?��`���>π	�`�*z	����9!��E#��[�M�-7�j|S�����{Z��u�d��I�����-q��}/��=J�'�,*�p�i�������x�o#�p��)����$O�����:%�,,7�s��<���(s�9��ݖY�6��d�E�_X��_���a�y2y���}����R"
D�eQW�,T�#��(��O�����H����_2���$*Kqg�I"=���Ż�_��KQ���)�2-���rD_�x�oZ��(�/7������s��3��y1�j�>Z���)'*�|N�ӵ=��{S�6�)������"D���o�J�>��%s��$�k�M�$��{EH�_c�]�Xɩ[����g���)1���ИDD�bl��g.���	g�d.i-&��t	�{�I!��w70&Ѭ�����%��9��.����ȑ4{G�nN�%٬>�����^��hXn����䘫���4)�7��$����I��%MR9�Q��zg'�IJ��%(*D`�X,�ĐUV"*�1�E�dP�:�hIi$EL��)��}�&���0�š��%��/n6����=��鞴��4�l͆����{;fD�����:M��V��T�nhN�����c�q��i4Lg�T���ё/���$��t�T*k�Oü�uh�hɯ��c�pcJ���=O	R-(RM6f���H�
#�0�