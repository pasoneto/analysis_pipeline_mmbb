BZh91AY&SY��6Y �߀@y���g߰����`㽍j  �G1� D�1�z�ڦ� Q� ��4� 5<�mIF� h    *������bA�&�d��@�5=4E 4z���@   i��&�&	��0`��$�LS2mT�P�h�Q���d��5�$��"� �<����I�%1��-��w�E�J��|񪪯)�D��#)D�RYD�S��m���
�wk@ " D�BH� 	"H���G���3Ѐpp��S��Nt��(4� @u&�=�B�0A+iژ1GQ�Q=��Ks����Bgn�l^z�):���1������#��!$j���!Y� 2ځJ���iA�,i��T6���[+a]�Z�a#� G��ey�]����gw���m��n[m����nC�ۖ%����m���6Z-��C���x����F�;��c�"w��s�ԉ�Pe�s��)��,[ �@�I$��z����(d�&�rdo5c2�[:�d<8�9�wI�����t��.�@줒Gk��^��ʏr5���S "��1��YB*�A�\��
�;�ȃ<��R�f�4�[l�J��6�]qmX��7rw���È Z;�4!fѵ����Y��q{@AӍ"A��h9V%mX�,�L���n�]q�/��5�~����I$�%ojV*������r;��6��MGr�wJ��q���&�9<�J��y��)%<��B�-TηP:��8j�R�2�:�s��I$�Dx�o�2o0�ڜm#q\b��u@=�w����ݺ�b�D��I%w��5��C���{#(���k�!O/P9�頄�����m��9���)�&���R6k��Af���N�SZ�v��d%�u�q�QQ�<M�I0�u�]Kα^:`=�:�|�_>]���_$���I:@�3/�f���2'q"ĺ�6H��Lw/�5Ì� w�4�1�i�F�m�����U�!;�Tį��!BrdJ�0Qr�(���*yX�aV*QE(��%�QR�(�E��!�����t�JV���J�D�B&d%K�b���M`R2� P�
�Ɂ�M�ěM���ԭG*������l��/Xy3��ׁ��^��Հ�T���� :��1��M@&C�B�M�
%!�����=�n�L�]b'y����s�G�g��a��t�"~�X}�=����f��q̩�KH�8w|T�������O�oV\�lM���� \��?��҅ĩ��v�D�jy�J�W{<��ϵ�:4.�Zq�Qh���_I���S�b���an2,T�k���~ݬ<ݬ�c��5�&̉J(T�R���}����In��#�iĪ5>�SA�o	��[���fn˄X����a�X��?�^�?���^S�b�,d��}|�÷Zv�ϱ1K�T䚾3���"`�8U%e&��;�I�k9T�'!�}��q�ׄ����El2q0�7ǲ���R^n�~��J&��_�n �P|ʁ!�Bf7�N����tT�QmJi-j�$�%�D�ĕg����*��s>��mMe�>g����5��)cS��O^'>u+%��;��m�Y�M��*j��(����g�D��J橕��di�R潈�U�yhel$����i�jp����X&��T�.-�E�%��9�z�L��m^���j�S-���Qh]G÷)��/:*�5.KD��Rc�m7P����C�G;FM|��>��G	�_��L��B�i�7�rE8P���6Y