BZh91AY&SY�c� �_�@yc���g߰����`	�.nu%<[` �9SA�eBIi�M45F���ڍ4z�����J��$�i=#L�� ���A�U<��U�F�4ɂbbi�!�!��jD	�~��4�  �0&&�	�&L�&	�����SL��M�����OH  4Ѧ�L ��T�F)8��O[��eL���Y�b��������㴂HJ��R!3!� �)���+�Zݤh��� @�4@ �h�  /u�U�ݔ��WVlWr��׋E4�,)�e�s��ȡ��7�:�A8��]������N�:ֵ9�[���ok�Y��(��E:�r�B��1�wp�c�%�ЯB�'&���c6�Jw�q<��>�>LS�ڜ5���;����^I1���)c�a�e����� H�~���0C���٪�o�:I�
뮺�R��[�wUU�����KL���˻��wV��DDn�owwkn�ݩ���0�h�z��9Èl{!��3�{3������bCFZc�_%S�"��������'��{��f#� ����\�����V��e.1�Z!�ц%����b�um0*ֱ�˳EE]��\f�@�j�KZ��3-3P�&y�C)L���8	1q���b!�5j��f%�R������s�qt�l^s���Kl�m���|#'�)+Fh���+��M0��Mᬚ���E�3������Gx7N����o d�J8�9��H�(I��S=��coAÓ�ݽuS38����G\K �E'�C	���^Q����1�~Nm̈nt�$ROg�LFr��%q�+��<4��1�BF'���HHK�U<�)�yOS#�����|�3J���
ma�b�9GZVC1��/��koE���u�<S�c6A��BBBKZ��*F/���y&�D��&`Qc�zVޝ�o��(Mn_OX�;�#�Ҷ칟HHHI� d�9�jڭ��9��7��y+]>�C��HQȘP�I/T$�u1w#�3R�����p$SDRu)�77�zt�q�w�f;��������V�y��%4��R��)c�u��Ү���h��Ց�+�v�k ���L��1$j�r��[������ɛN\��j���U�v�j��nZ����}&�WX�ă�%��s��2�m�<5ҷ6������UJR�^z�D����g]yF��|Eܢ���%�H �A��((F!�	@\��b�lp�Y/{���פX��.U������F����u6)0��T׺���C2I���s�����Ϝ���u<؜�7};��]{�c�q�ؐ���Ij�W��Q����ˀ��wQ�7泇��=*|����j����ޢD왞�qс��y�<�'�VL$�v'p��U˽OK����X��SXR�^i�)����w�A"�ɟ��6��O�'
Y�Ւ#%9��m�8���	a�x��v]k9��T�Z���ot�q��T�@�T�x�@�{8J����R�Vi���ã�ɢ<��3͙$���AR��ş{bQ�f�[�<�s_���M�it���l��l�����0��(�.�X$��ӌ�J�q3-d�M&EPHɎ\��·�p1�Cktl���x58�%����?�����|�'
M���������]�^��cEk2tRs��O�-�&/k~-�$�;,9�0L��~R��y�kԲ�OZ��Z�k1�S�F��-j����`*ο����%U�9'�]<�t�,���ϫc���,��{>\'-�Ζr����i}�,�nܚ0I�eڎ�R�I�p�΃(�b�Ŋ,X��QE�QUUUUEY 
��06 h�L����:XMt��Iޜ��2rj,��'�:u�\)�P6`NV��[J�ԁ!Trb`]%3���$Rrb��,�Y3p2d�U8�5eC��E";�ֆڃ�Ġ^�f�H��1˻Q*<N�~�]�2��J����?�w$S�	�>
 