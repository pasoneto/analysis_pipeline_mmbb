BZh91AY&SY��B x߀`y���g߰����`�y�{�GP��T�$�S2M���!�=OS�z�=OQ�i������~DƔ��       "���5@2   h4 �AI�ڞ�  h�   9�&& &#4���d�#��hB����z������z&�(xTgB@8� ̔�s ���[�`�ّX��%)LɆ�m��Q!
��I\f�K���:��G�6�/ޱy��@P��D� IAJP   �j�颔Y*�q(�b�+Ń	��A6$�	��;�le)r�4B�A���Q%�PS�dS�xr��DRd���)�l�>�t����I��M��2�X���2�$ +-�P#5'0���[Lg%���w8�S$�)�D&I%
�ZH"H�H$��$�D��I$�I2IXJ.s���۷�!	��������Q�8x�xw-�x[���}���/���� �J{H@XJ$J˺�
Fb�1�	��T1�.�ul�i�{ղ,A��@o	%06I�GfJib�	a�\А�1Z�-��(gki�g,��fS�ᆓK�Q�KE�ygr8 �[Y�U]�1�Ԁ�3q��-�$�K� m2lsI��!�4p�0h�7,�\�H��i0na6������#��槢	$�,� /�p�UIX��Q-$Ӽ�z�k���b�g��L_'S�jl^f�;��I$�I5�~2-o����/[�q�k[�qmv���-,��rI$�z9��-�ݸ�Ylj\T5{mkD2S�LI�����,�6�R��a2	�@�����j7�q�ͧ�q!m1΢3#,���.�H ����4�;S��p�<ڽ^�B:�Bx�����i&F��NY 5+a���/����T��ѧJ��N�i	��p  Q�4��Tw��ƥѦ�C;�G��3����&���7X�A�$�&��z���~�I�<{㲐@�ēt�U0`��0k� ��4����B`��0`��6S!00����	�	C�(#d!�L�a�2���5V��8� C`�lZ��4���������yvq�X��wS�� q<�<͒���a*��8��K�W�f��) {�aА��\��z�v;6Ș~G�Ni!�rh��z��4π[ p�N�!��8�^��!�+�_0�X!y9`\
>1�B�Z�ӆA��%a
G �K��}� 1�xV|&"Z�ǳ¹���(	j�%ʚI51�(Ml�� ����4G��dX�B!0�� �y}P�5.wо���M
(j��H�7j?��{��ޠB��ȳ�M�)��j� �s	�W�VǦ�i�p�T�.�T58����^�B�7���ܪ<������MUZHK�Ba����$얷U5c�#f���X�T���QJ ��ROOD{�
VD�7��-۞�MW&v�FdD4X<�T�%@��.�P&gVX����W�����{h&��Ia�r@2[׹�(�L�MTu8C���=c�(BBb ^0ɓ,ŻK���T�L��?"�.���ie���H溄�!�aV:�*k��!B@�p͐�����-�:�B���Z��嶌�ѩF�,�Ï#�Pپ��PB�A����LBt+�^�bJdR!���\�ف�T�+9fu���
b���ܑN$�y��