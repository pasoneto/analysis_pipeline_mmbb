BZh91AY&SYҐ67 �߀Py���g߰����`���v� Mr   ���?T�57�m'�02hz�����R%       9�&& &#4���d�#��&��j��G꘍  @  挘� ���F	� �D&�&�#4L���OSCCF�hM4�UQ��t%@1��D��0S��(� Y�J�3t��"$<J���Ɂ��|$���]�R�������c�Ɔ�y�8
I$��⍵$�G	$�H�#�r1�q�W��0��	8�f���!l� �I�[̶ض��]���W�������5&𨙛���S-����maD�wUy�U���wwRAzc�q�0�H=�s��0����I%�6l�Cd쥍z5�w	�ah� e����R�����)��g�I��| �3zR�Tk cU{%qS��j�Q���@�KE� �(*"�o�	������T��b�}xx,��n�3��fݯ��sLI�z�ח�'��Pet*g�T�3p��N&���"����]@��jЕ�C0��0�z�X&4*^DljD�`�eg��'Zd�va��e4̜��5���CX!��2#8��`5������wCxm��wm���ۭN(5L��1h�2b�GO��7�=��J���Xf4m-ט��9A� �z�Ò8 ��]0v���C�w�W�،W"4��N����+���8$n1�+�~g)8������CE�9�j���/4��#[=�(�!�=&��g�"GY	7`�Y�f�5�i�ل�V�Ӈ�A���(i⫨�{aeq��K��
UQ�!rᡞHk(�,R*��$����C�3fj�&J�轉e���Ȏ����ʄ��=�{n3v�.�ԗ59�ƹ��@׀�sh�n�mͲ{qX��M期:�[�t��{�s��'�A�D�H ��$��;G�B���)4~�N��I0(R�-b<`)
�&Ef1�)�����$J�!�6T)� I�����(\��!��c��P� T	�������t;�q�b�z>7	Y�O����Ȏ$P�?+�������^�F�X�%�by�x���m(x$�05�G�r?3Q��hv���Jb�t"?P�ᾗ�A^�F�|�8�D$���Aʡ�ݻ�"?A���I����;J��ИD@D�;J�|2�I<Lr9,H�����;��R'��i�z���5P)�
$4��K���	/�'GM	��q
�s�0(C0D�/��L��)��BF|lC����� X'�5쇷�%�U�$���!�LQy΢�0���C����$�w䰘�.�;�<�Ϥ<� Y�B��re�xa�f�F��� "��68���Gx�t�G�=@}����;,�#:[���(��b�����M�¢�b@ӦZ�ڟ_OPd�����1��Pp��4�!� '"1"a0PXTejIì�sxnV"jr�G���;4.H�C�k2_I���:�:�*��jw�C��sȲ}�SW1�@Q�)�yM�#�=5KIm���X���������Zh��N⓺M��=��C���.�4�+�yJᣙ�Dnq��j�3'��X�YyZ��&+c�m,��D>����k(=l�������)c=�!/���Bmk����:?�w$S�	)cp