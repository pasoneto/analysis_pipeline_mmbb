BZh91AY&SY�W�� 8_�Py���g߰����`�|��˳(
�|���HPSԙ=L��4    �� ���J� d2a ����B)�ꪃ�  4�     	L�E4� ��`�i� ��4��i�S����h��i�@"B&FSѤ&2�S��!�M�h6�'��!h$i!c���Ő+DX$�:����� B�(֪0@Z��QWS%U�)F���@���f5�,��w*��BI��U	( jɠ   �UD  ��ӻ}g[yH�l����g΋_%c��X**�(ޝ�RZ�M*��1^Sd�L�L��
�����z��Ut^C�ӂ�Q��D�������a�v�!k��X�r��Ah�߄2���lE���6��j^ka�b*)��\����~�����y����$�T����Wwwu�X_332��]����U������uT*�]������9��i�k�vvr9�D�@!|�z|=pw?�J`�(ߣh9�Y]��難��Uk�uI�t�5:5G��MF���cO&���M���8qGEm��G�FDBlm��qR�Pp���-뼑U��2�	Q%�E�g�ADb(�傖YP50�
��Q4TU�yf9��m��yo�����d#����m�)K����4e�ib���F,��2�[]�*�"ȉM$Ã"���t�� ��w|f�������A�Aի���Զ�m��y��N'�b�CS�2:j,��bPM�[�pk���:�g�
ffffig�%�T5��.#�ū�D�`�����U���,�����&:t�D�]EL�O��� m��!V@�.���k���&ff`��'�\��隲d��RYJ�OU��l��aԗ%'V�m��+<�ql�������ə��s���Zu��9�H�1c�q�j�/�٘�Xo��t =m̩�<Wj�k,*[{|=`vm��:�+hƄ8�ǰmH���#��;v�������!�	�	xI	@""�<����\jv��b�{~e�2\�Xh�Ʃ0�9vYk5b,���͗QEJTT�S*�e]YQEET�TQQE"��Uc��D�&d$���E	J"0�Ց"3
d�b�F�6wUx%
�J��U�
:p���ʛ�;�eroo�E@?���]f��P��Ӥ,�.xPG@ab���d��k p9��`\q��2U!��6�1�3��?��9'T�$Oih�Ka�iڦ_;o ����jS�&n��d���3j����5lM����&���5��ڊUR\��Mdy��ÏDc'r��	��_1{�W��GXȠ�c��ʋ���>I��¦Hj$�T
1|�,��y��K��?+��&�4]�h�/�)RB�U�f�Qg;��(�St��tE�7�B�3/�7���?��5��T�&'9q�u�l|=�gZa�6�mɠc}��84��`|�!��{���vS��Tk4;�	Z���w��jςw�Ӎ �$���"�tW���;�~rku���bQ7:��9������nL����|<��[��`�\QM���/$�wm����O�E�)�]Ԛ'�3���B��Xu��>��*���D�'TܛP���+Q��g*Y9�\z�s8�Z�����S�s���s��ߴk�!%M��y�O����� ��,44��PmM���D�j<4�T4�IEl8�_�N��F_45��p婶���2�SN�QTlu����JԻ��4��M�ܫ9���kω����c4�r*��g��7�z�OZ�y��z�'6�=Ƈ/K����Ε-?Mn�Q:�
{u?�w$S�	�z��