BZh91AY&SY�B�� 	�߀Py����߰����`����k�R�P  ��� ��I�ySI��zM M�   ��jS�2��&����E=�ULF�& CL 	������CL� �C  �b@ ��� i�e4@@�@4bhaBx�I��F���zHd� ��!���".'} I*�i�!Q��@�A`U��
������ĲX��s`qQ�P5m�%*h�@B(�} �1Hx�×w��9:L�V��Z�8 �@!� 0 �@ 0;�3�$�$��$���'���ˊ�z���Zx>��8��V�����р���SLy���V�/X�ޒ[ͨˇvlD�L3��-�[�h�=�C�H��_oW�.��3�gk�Z���Q�q���w�4a�랠�z?�瞦|s�~���2tL��W0��L4�ż]��!MʺtCD�B�U�C���7jٖ$�f����F���{$�[$���� �{�ae�i�z��3ٷu���Z������w��332�.�32Y��fc��~R�DN!ᨈ��D�$!�gww��N��;��"�;�`�!��m?J0��٦������@��?�S�{G=k�Ι�,y������T���s2�bdUK��s,Q�X�,���v9�CzD�^���Q��8ÎQJ%D�dhh[���s-M��		�Y2�E���� d(Bwb��b ����`�$���:�f�*�%����ɹ��a���k�<� +-?�(��%��z�HKI;wM�w�b�Bj�(,@��@�̣�ܠ���Bٕ�lB ���0pC�6 $��ȅ�0�E�Q7"t�z�l\�J	�Ԓp��
 �q�������f9�f�rJKN@�0 ��(sy=hs�6�t�S��30ux���$���%g<��A�"�`�q�8�WB�ᚱ�8�B$���'9�!�N�6�����+j-t�'�Y��C�z��
�I/�����5#�6x��H��l��=0b�9)lFj�lr��	6QC�;��On33DTR{�;i$��$�1afQe�I�Z�����.���ถ͘Q��,C���������,�Z@�0ܨ)�2t+I$��(�@�`�,a�aG5�.;�d�`la�tQ.�8���)f�`�vt$�Z�㤒W�$��l$��kg{K ���q����,D�#	�!�,��f�����$� r�q���(80�) B3�s���)8A��G�mv��6�}>G� B��P�d���S��OJC3�(�j�z�%��,efوތ�TְXeA�����"A� �PRTHP�	KEn@��f@.\(((X�Yk�ЫD�"X�D5cg&��`b>[I�b�3 3$3&d��{��M���9�?��z��Fj�w�E./yz�B��WBB$�Un�8��Wk_0J�5	�$��%BE�I"�1ba���|�.�*L�<IQ!̇��H�_)�7��`�>�R�����ą��7r��)��24����n���C�*?�39��v����(S�s�_�7)#)�ros5>�cM;�u�2�x���	����p���x�o��n,����EC�
W!
�AG�� Q��>�<8�����u���� H!"$c+��v��ښ.oPV֬�vtaP7;��B��+%�?XӴc���f:2�Tl�
M
	a;��~_r��Js�0��z�x��O��;�h���a��`c�����ϙ�N�Q��� ̃�?3xdO{�2S�;�����j�9N����Յ������?3�.>
}y978�>�q��*���~�.ae
=L`�4�PCkS�����@]�cB?9�R5Qr�& V��$�k���H�Wg@�)i�P� �Y��>����R�7󣧍X��ì�<@���%{�@�n���ޤ�Y�s��6@                        BI�&D�դ�%+IJF:\�8�4Sjx8S}�D���1iۨX��m����,�����7���=��pt�s�|�.1|���B��ԧ7�
*��r�p�0)�A`;�ttGBC���a�<����u@#�4�Z ��
U�,�)+��TL>2�Fa������,��5�ܑN$5гt 