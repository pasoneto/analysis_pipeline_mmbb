BZh91AY&SY���� �_�@y���g߰����`�{ܒ��U�P ��D�zd�������4��=A�T���      ����@ 3P  44  6�$�      �bdɣ	�bi�L#0	Ц��F	���CA�#F�%���`�@ ���. K2�WʡB?�$T�4%$�&`��i���&���#$�V���a&���=!�v��NuW�  �@D�P ��� @"�mw�(�W%q(�b�*���膱ID�ʉ	�^�jR�gjC��כl�z��a�	����h�")��0�\'JnnO�ټ�}��	�L�/��$g�C8�0�:w%��d�$ )-z F*G(����8��_9  �` �`��0   ;��    y^s��Y��`���ϗ�>RnA�2᧯d������[�թ(����S���a6�m�-'iۉ/!"���1-fQ��ͨ���Z7x�ܰ'iF1�P�![0%�َxP;�ہ ���J]��u|�,5�P$�L2�%n;\��j��zil�rh��ůL-I^8�'V�5'K@�`�uBF��Ɖ
��o��b:�$�p�u)\hU��\F�=4���\*5�M*ȶt�6&�ˣI�Yq��^g(E0o���;d�.�3p  {�kw[J��S��W�oT5��Ů�{��u�%
7�ם,�T/�� ��6�x3�P�����CZU����R�OJ�t��x����� ��ڕ���&8-�kq�i���m��^aZU]ԶB�+�|b��,��  Z�:�W�Y�b�U�����),��M+UUä�divm��+2���Z���-z]4��R�#%S�X��t��Mo�n�5M�v^J���%�f�_H������UܩUj�J\1&�/S���UUWL��l�Sd����L���&�teJ�1�߼<F�ߩ�ؚzhv�v((J$x�G\��ʤ�X
&Y�40a��40`���*�C	�Z�i�V����j��Ja�A%4��  F�!w9�B�]�[�i	bC).`��_kl���拣�r�;T�-~�|U"�D�.��gZ5R<��j�p.��(���1�%�r����R��,��%�SXW	q{����HB�P���^�?Y�b9�.�� �<��;F j��"Ą+т���Q�j婢�:g���!�h��l��dy\�HB��Ak_s��gU�^��q&�/���%�d�f�9@��j�&���D�-�Nby#��`W�$Bi i�� q��G Y�;Is�3��YP�)	��4:�|:�����@4�)�
Ð�Γ�_�[�n\
�a0��73�U���9���&�ȿ�馸��)6���h�<Mm-%�6�4���]g�&1�H�ZQSRC'5�{*T��ii�&�% e琧#�ݪ�?¢���cȆ��
�c��T���Qq�PQ$�	LG���PM��zBa�d%Q&��� �[i�����a���鎡Ԏ5.|��<�"��S[2А�p:4�\�IȐ��.�0
���ett
�� TmT�G-�%h�y-�|�n�O��[��¹�'P&�I�.eT�+��D86��3`�*j�$.#~˅���m� �Rb'����(]
�ʚ)"<��^[���N������g���"�(HF��m�