BZh91AY&SY,�8� �_�@y���g߰����`��GL���		R��M54��٢��S����=	�OP�ѣ�56�Ғ��i� F� � A�~���4�� �!��� 4�M6�OԀM     �bdɣ	�bi�L#0	M2LI�m4��'� hhڞ��H%Ԓ@1!� 
���� J����3
��		�a���py%�i+�h,��|��|i�L���̥ P &  DA % �үCM<����9?q���^�6!3,j�I�ɡB��}��8� ���Xa,$X׶O"(4X�3`���c� ��6�����w�?�k�Xՙ���$׬���x$��L�ZZ��L��
�g�poz������>x;�3�I+I%32�V�IJIBI(����t�I$�I'wuĒ	$�I$�uQ����!2`a�ㆍ!����;C�n{ u��x0�<��TX~0�ffb��ew���h�CS��&b^S��^Ijf�%yG`9�� �%�""���j�)|�ӮE,u���@�MQW�2�uh���d8T�e�d��J�	�����K0g��K@Y��J	$�*B@��3 PȖ,$X&vQ��8T�s" �$�7:D��J¢��AE���S i�(M�����#��II<{Y�=WW1�{AL���'u	�3)�s��lI��,D�I$ڑ���*_N�Qjr�"[��
i�])Ǒ*��c*U���I$����v�����׮��j�]é3l�+p��Cf�'.dф'q�PI$�I�<h��̶д2t���mE�P+�e���x�F��I,Y��]�UV����lL���w
����~�vD�Ȋ�ޜ˪��آ�Y$�3H�s:Z��
b�lu-����a�Jwt ��mV]l@Rє����Ž�ck�-˪.�f��B�-bi��s:��x.w������X3Llc~��bi$( ��^栩1'��Gu �͉&�U0`��0�0i�0vb!0a�h`��C�T`9��$a0�aZP%8b��D���"^#)HCUk�e�BM��l lU�0���~�#��%��Zk����P��[���֨�������>T=I�I����ȹm�~@k:-:L����	J�a���ʺ��P��������8�E�����Uh��bbd����c�)�)bs!!oD��T\|.*��5",�!�W���dyby�R8�^����z0Us0m%���U��++��!�	���ܔ&���8�a��I��u���y�Qk�$Bh�� 㤿�*z��}`fa�6�7).*����QC���Vv�P	
M���ZOa�w,�d�'�A0F	c]���T�W� �%���TeP^��1Is04C~uQ֝�1[���$.g�L�q;I;��*��X�Hř+��ԩ�����(��`e�"���r�x�y��: �~A����F`D4X>��(E pr�p�p&g�z�abfT�_㞳 u�H�8�KW<	^4G�M����Zq8�7�%�*$����Mp:}��	�^���UWG"�- N3,�,N�^d2jT��N`�݇eb�`��ᡅ��)`(��^ud$+�ue����h5����r�S�l�S�1�3+LQJب�"S+�x�ve�R��с�bb0�����)�f��p