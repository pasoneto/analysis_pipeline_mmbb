BZh91AY&SY,0s �߀Py���g߰����`
��﯍|��� z����!��	"&��F�Q�iOQ� 4� 5<�)Q�       �<�Th	�bc@�4�a0M2d0�ME4��h�     �*b��@4� �h��P �$	��mJ`��=S2!�4d ��4z�]�qj�!*���Z��%QnT��ǘ�?Q�c�* X��}�L��WS0 ���E/�P峦���&+�3�V  @ vwt�T����*���n��n�����@  �f�0(T��hRu��Ī�Ou)2� 5 �y��t��w��|�]�M5&��d�l/���a
6HE���3r��&!&s��5���#F\~�Ƈ��}�rFx�N����hWn|�F��c��b��M�w�v9S�T]KEu�g���JvV��iE�y�����\�)Q�Ym�:c�e|�R�ؐ,Qv��'��]�8_�U�Zֵ�fff�< �www<�����pY��ٙ��R��b"Bf��֯#~�@	00�nn����$� �2��aӞ��yA6bZ��JL��y̦{rvb�30�Z8c6q;kaD�-k|8�]>�Q/<}���ٹ�5�v�&�g�G0�L�eX45֫i[��5v�w�"�,��P��vb��͢.��h%�t�`m"���sl�����4'M��]��|���S����8e<L� cp �S�8$5~t��p	px�׈ �������O-ת!x	�F<-�jњ]�ՎU%�p56n�JL��6qb�@-L$�kr �kd��@�,x0�l�\J�m�`��{��f��FCo2����P��m��vf���I&s;T�z��>���C؃Ns"v�,��6�n���9H�!!�S	�"M�ôe�(���j@�����k	�ݣ�ˢ"��Q�w0I$��a����}v'�/���|�ᶃf;r��
����M5_]���w�ܻ�_d.�;��g�!�n;v���$�\z;�DX#Y���h��y�m9X���܋�0��%�li�/Y9�k1Ɨ�x[uv���J�&��IL�R$�C�3%����`��v��b�",V׈�5���y1j����	�7/��R&�a�	���!�ʡ�Er�rI%dc�.	��(��1�u�
�M�T˶���U6��ݓ������he�l;�=!P���S!/&K��0d���xI'��9�����ǵ�(�I��ӧ��^�Z�E��VD��)�"�^k�K����g�2gEMїʖ���P��!�[���˪������*o��x��:��{㼁=�r��4�z=��\n��:��DE��J*v�va�ǓEJ{�J<�Q,dX�"��^1!3	a�hH�7P��@P�Q"4X)Pi�-��ID���ZU����Fe�%�j!u�4��9�����"2$���c�y���Sʴ��x��s�������=�}~�i V�q:�������e�*=� vu>ih��,�G�w!�}g�fq!��� /��m4�_��O���ED{����>rz͜ԤlORJ���o�1�,�0�/��a���7G,��n8)�4
	��J�Y%5����Î\N�e���3�n"-�5���\M��c��4~ݷ�=��>Q�T:�
��E����ǒ��h��.�:����J��:�9��@J�"`��rT b�����i��Ptj:�m�X㭬�}�)i�~҂ -���i�n;���8����|�",B���}K�;W���.�LVL�o�n���f �38Hq<����st����; �p�c�,u��5�3p8�	�n�!݁�q�(h���r�M�V>^�)Gyx��(#eOȫ��ѭDu��� '��f��EV�bK����%ht /`XN�h����a�}�CCbP�t������͏�C�yi=�Ks�Y4�&�:Pc�w��
�*�����**������UEEb*(��U����*(�(��UUEQUb(�QQUUE�N,�@��1�9��8��ˍ@BG%z&��!�Mz�I�9Ƶgw�VH��n����t��]�� ` ����6^�R����w���O�����o:Ir�̽JG�#w�ڜ�a�j��[�l����t���	�)�U��w��U����)�a���