BZh91AY&SY�� �_�Py����߰����`.8]"J�)�TAF	ݘE"h04���&�=G�0����=O)�%O!H�*=F ɠ2�  ���M  H�     4�UH44 4@�    ���a2dɑ��4�# C TI��O��G� j ���"|��!��q$��'��i	7����{�\I��8�#�&Љ�<ĥQ�T�0�ZB��BH����ٍ{"�,Կ�v���A *��I *�B$�
�kP"uoܥ.F�&�FR�ST�(�|;:����k��.�+���V�T�Ӭ^��4�Q.�nw�\���CNh�8�vѾNl|�D�2;�1{�x������(^����ǩ׶�O��ߦ��������5��Jt�!)Pq��ʆ�4B�bڨ�D�:R*�I�|u��S3�di�tp�"�|��߰��U��Zѭw�wߓg�4W�������ۗn���f=37������32"79qy��Y�̬31���W*���3"�]�y��-�/�����@F����8��t8޸��j�k���ECr�U$í1C�W�>�I$�D���3����}�_�d�N�ڕ���N[9�M(甤�T�n8#Q�gF�1	H�'��Z5�jθ�(���Q�-k¦���ʞ&�������l��2*�����Һ�ݛ�x��~]mnǢ���;)�^���[�n�'&�7z3����]K����ot�'��S��Ưm��,g���h�$d����
,��v*�ݍ��M(�M��S�V�y�dr�٩ӆb�cy�`�<`2V_f�Dx��L̓g����m���y;�p���ӆ�6�r�͚r���0��Φ�،(���QF�,�d#����[,��\��T��xt�vESm��[�Iٲ�$�8Q�5؋8x8`���Y�K6I��6A�$F�I�����>O'���/�oY9���0�W�m��r}�2Dp~���Y��$8p���Qb��2D
������,�QF� d��8e�.MÞ�_U��!����nwO�_X�m��/�Dj�0م��,��3
�(�Å��KTA��n���4��a��w'M�[�Zq�_U33T.6�MtQ$�l	0ل:���3�D�^
�0�W,�Ԭ::
����G��I)��c�x<Q#$�F!k��Yl蔔�V���:y1����;7:w�-�ZnZ�l�^6��e�C!B�8�C��@���$��ta��a�  ��u�̵-D�,�IW��R"!WT�R�Xd�n�d�Y'?$���O���ǳ�q��4��E��f�E0��0YRR�`�J)E*R�T�V2b�bp�͌�YS	�h�jɚ��Zѡ���i#�*�+g7����(�l���\`:�K;>�|�m~��f��Q�G���^&��>Z�>1A�A�&��۟J���_�i#O"y~��$��\t�����/2 ���q����/3p�OY��g!T�d$C!��;�*�0�!��X&�d��t�zq�xk��v ��P)��!A�s��'}R�ݟO��Ն2OSnd�ݫ��v}}��9K,��3WqjЊ�虤�������I���!�ԁ�TB�g��,���\+"��{�����(8�����V� %-�
QeU�aϷ�B|Q���ߝ��w��	�g��)�V'p���3�B_��=�k�qϮ0����æ]!�s���+g�9m(��e�BP��vA�S�9,p�
=+R�#$�/�wY��rA���V�v�n��b��A]h#�t� j�H�7�ED��D��K�XM \�7p�С� hg���DAaIc)�~�Z��#�n��:ђ�2�̛���r��$ߥ�"�qr�s��-�d�$sxm��"[$���7� }��İ?d�1Y�f���@�#3���X:Q�%d|�v�9��T��b��V&��T�U��/O�`                      *V�ك'�A�P`��(6-��*\K@�،�y253B�T���r�#k�e���t�9ua��g;,¸kU���y�Ʒ�ѮƽMwZ��ǲ8�y��,����i=�:WCwĵ�P/(���J���3.x=�OЃ���q�IC���<�A	�����y �HW��?���)��`��