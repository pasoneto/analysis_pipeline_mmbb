BZh91AY&SY[�[ �_�Py���g߰����`
�}{��}=��  �J��*����=C#=O(�= h �� ��BI4h2d�    ���  �     )�(5	�@      D�)�4ЏBM20 24i�jEd LiFM<RzOҚ=O҆�4�����;�����BUQ/<�� ¿��T�>�`��^E� T�"p.\X�@�.�� �+���)m��@ A�  �wm�䥐�Ad���$�ܗv]�� A��|�6������V#��R(`"�DL��[ă~�j�c�U�$�ū8���ӳ:�!��z�����j!���Ԩ���1�y��2V��?d�	o�>����;�O��A�^�O|�^�P>�.�T�R�}��w����bȷs�fQ�z�w2�a�"�QNgT8�>�űc�M]��_8�P� T�G�$�!VD|��Hw�ckWE�n)A%(�������$RJ�{F��ԋ3�I,ř���wwv�{���� f bq�n��oDP9áۙ{�d[���]b*R�9)����K�f*E�4�.Y�Ao���C�Χi@��U�W�E������h+���5[+h���E(Y��wad����j�	�.1���q�k
�J �hp���K�^���[�K4�d�~R�F�j:B8]��Ya�hn���k�i�L�5ts6�04l�͢RM�V�\��
nFCJ��ޘ���c� l��ܯn�7ۨ�&Z�Y�Z�L3�s�s�]����s
ĭ,���%����A�� 8��h�E��H���3^���Ȣ�p�.͆�:��$O;.��FN'2|�`)��^<o�z�����I�]@�z�����X�ֵO���s(fn�Ueߝb��^B�ӡ�[�
������*~��Ot}�=�0�C���Y�����x��I7]m}�f\�˯�E���ۈ"����A����^a����Q'1���g�Q�5$M���՟0�f�%S~=rI%1օ�J�.�"�e.�	��F�O]�z-�o'8z�5�"!��p�~�=un<�ۼ�c�[E�;��ɎY����@^�PI$w{}��'#\�t\��$f��G	�+5�0�����3�yb.3B1s]v�����q3p�r0�D�I{9�fa1�����8Wl���[VX����{������G�����2d�����b:�:��pC��5u�%te�>Ēc���%��d��&�Ȃ�ޞ�-�;۰���/9�Έ9۸�b�%�l��ݲ�cO�����y�ڨދH�\槻��$T�X��'^h���T��.�r�хR�C�N��*v;����A�!I�,YDx�=c���h���۸C��6BkUA����XF�ł�$L��
$X�c�Aj�(�q,�PRPMF�� d����ue6	q�R��99@�I,Hg�"����y��T�!�8۷{��N�X����*I��&Pu��nOϗ���h��ׁc�W\Vm>ә���o ���.��1�e�9g��V���*#ޔ���q���2�ٸv�Qp�;���!�P��� _�_��8����
>��;[�d�*�`	$v\^=��$���2� "B8ߎk���z��=�W���?��zH*&F
1�fRX}J���!���w˽�qz��N��ɸ(S0	 �$A#V��*�ԗ��A=g54��T��9�����&è�s*=�G��`���B �����g}}����*��vB_Qjn����Yå2
��r�,i7&?����p������#Kb=7�Ð��Ur ^õlu�R���=L���H��;׾ŋ�a#'E5�[�E�4q������<
�=X$��ɸ}9�G8�Y�Cf��j���p�t�mV"r7 /hP��@�Ù��?鑠d9IǲCpT�.����v�Oq��՜pK�*�eQ�)��#�w����*Ҫ�*��*�*�"�������+J*���*��(��*�*�@����J*Ҋ��������UPV*�)4�릂ÊzJ�{�@� 0P��Š�����cA\gúB�t>��N��	P:8��yк�A[�H�rKj5� $jh�kA���w؂ �T3U�w�j�0�!���t`k���#qyG�S" ��݇f��E6��"�H�
{K`@