BZh91AY&SYp�N� 7߀@y���g߰����`	��gwˎ�  ;�>�h���B�F��	��4��� ��F�      *=��&�41 4��  	4�	LQ���b4z�0@�4S�SM(y��6��Pz�  ���T�4M�OPM�bz� �����/d	 �PT
��!Ah�&{�$f���	��{��tU}�H�8*&���H�RYDʍ)����4�T��_ P �    ����331s.
�*�Vҭ�kU��^�ϰa�N��ܟ�����x���+� $Қk%�`eB�	��`�Ծ)�)2KF{m�w�]ޕR���tͦɯy�#b�O�PJ�(�����Vi��^S4���UUUy˻�M^K��]����a<8�
kd�Ծ�哲]�Sn %��\�nBN���<>�:������o6���]uUW[l7�\�WM���U]��t��cd5��.�~����	�"?O�N��;>�\�D�/Lx@�j����t�9�(���P�H���y��8�n�:Yt� Z��%��#`�R$f$�j�B^��ҍ�A�7R�a|��ZJ��3��#Z�	X�$�wP�"��LdFj�U<�A�)���0V�ruK�J��mf��o|0D��E���i�댈&0*��[�l��4��UP#�*��k^�	�s���k����t�.���':2J�,َ�"z��z�N�h�<B�w��;��"2S�H�$�$D�-D�@�S�mV���=�p��ø7i��_ 2׿%:�$ G�^�Pӵ#Tek�nsV��ε����@=;
}BC�D�zuW8��H邈�|ר�D���D���(�a(E�
V��G����k�T���B�%tUz���8��=�>��i�a��33B	PrļZ��I�nq����/�d�K���#yC�8�i�0��7O�`��-Kk��v���/Г�Ͳ�m*Dj�+v�v9��b-f��f���¤�/Nt2�e�(,��n��D|Jx��qx�*i��qٙ�ͅk����?X���QJR�W�UP$%,�5�������̸΢��C�T�;���T�!&�H�%68(�H�d32`5!,&fɍ�0̀p���3Y���!�:���c$�(�9�m��x/��\�o�5����[��- \0sO��� B�\���+Ɂˢ���R�
�Ϗ��n�g��v,�`���Qs �y�����zo��:�`��d
��"E��g��)����W�L"ZG����$lD�� Q�ZbW �t��@Mfc�?5�	2X`5��t_&x��rf!%Y+��zkϒsfb�Zq�Qh��辩�ʦ$C�QU��"�O8F�2Qe�M]�yxb�#�މ�\���R��D(�&{�uF�3��xݲ7M~`�e���a
jFE������O���`�{	 Q��!*D�3�y����W�嘤�'*��N�í<�֘�ӽ9&���~-iȑ0i8U%e�yu_�$��R$�I��#�u9�Vn�������P�`x�����%��7�LRB]bl�b3�/_Y��3bj�E	�W�.�7�oC�5�gxB�8�d�)�K�&U�N����V�$OI��S{a�5��#�����湡a��?n'B][������q�+$��9���SID$%��;��'`��g���,X�2��`�F
�bʒTUT�J�N�s@�*g��F��.��R2�F!ռ�2�QW�L�(v�v|0B��^�j��R��9JWgQ�"g7����VZr�mnQ7%��q70,橩2��N�ڙ�)t��M�*i��w3���d���X��$��W�c��M�����q�rE8P�p�N�