BZh91AY&SY3��� Z_�@y���g߰����`	_z��{  � 4E�D���O�����2��� M % I� 2�    �����  2     MHD�	���G� �Ѡ�bdɣ	�bi�L#0I#A�L��`�6I�6���jzOS�݁wBB�"1�A�|��&2-��#,~�*!��uW�]$NJ��Dg*$�u%�L�֞��d#��8�02��� ��¨��� � �   �
�̀8�û�2���3�qi?gO�_R���(�־����o0.p(�I,�F2Mcq�^8�(�cK��}��ڪV�<n�o�9�U;���i�^Wn���wwwuX�[��Y{U��ȍ�g2�f��v%]����3�Tb�IecGI��<��z*vt@&�S{d���\��NmX�ت�]�\VYY]ڶY����j�����<UUNp��UV��j��T�����mۺoBB0H�w��Ş�G+*d��8�	���0��HǞ3����2:�oj���b3�d�8�^�� �!R<�W�w ��y\}��<��@u*��BT�`�<�Pq	C�\d4
�3��Լ�d6BDw�mA�ͻ�ax�҉�H���#s:�f�g��F�è����G�*,bp��8��.Z�x��4���m�8Y���C�A˖�B�1]h!�iHA|���2����׈q�S�bJ��"��z�^�fQ
	�GR �r�9�һ�0=����!Ż��8��Cx-
ԅ�\y ͑z��Д(7����A��à���Bg�[�B8��U���KdGv!�{L�,�ް�z��z������؎_8�-.du��<���k�y�i����gzY��6h�O��l�B�ݡY&���r����}��LU�pc9�P����љ$�f�Br�$7A�Cd�	F���Z@Ș�����AeG��b�k���K��̚��Pj�p���	AC���2�3�{|�����6A�.��i}KC�rs�:^�ha�R��	ۊ���UTJ*w�9mC3�(ĵX>�J8�T��ȴ�d�1&l��	ip� �R�Vc�#{������ �%R@�-kb�Y*R&���J%H���w�!�$�3 ��:{�#���#G����Z�����(�^ʽ=�"���J�ۂ���x�xYf��Kl�r���S��,�����5L�]�H������������St�H��H���|Z������{��D������)�����ĉ��l�A��4���Ó�����"�ʔ���FT��5hp��D{%���Bzń��b:�!��8�,�ʐ'�DI���-�"�OT�(�妟<�b��?\�.n�D��T��	E��ɤ�I�ط{�#���s-G�SDd[)��-����KC���D���Z2Z��͂��_����ڼ��頤��N�=�ϰ�ޞ��y�&)t�;_�yߛrt�St�T��}fJ�=g4�kD�nvD��{�H�^����aGU��[̛�%&y��)/6ë�b.�7��3�>���Ė~l���E4��ʸL�����3�B�5F�2'ޗ���U����|9�U�t��"h�K�)�u�`�a�>��O��5�t�����uq;]�
{)�d�{癉�����C�!�8N�韨��PPPPPA�#D
(,X�bŉDQ���c��H�S<�25�u��#)Tb��P�I��Py��*�g�(#]����G	����c���(�3�F��ږ��e�bl�ZQ�Xzr�����T乫FD�'�]%�j5�O��c:�t�d���c��zTr����yʑ�(RM7����H�
s0��