BZh91AY&SYW5� k߀@y���g߰����`z��N� ҙ4e�ID�E<)連�z�h4@� �M�4��h�2�  � ������        ���Sҙ �M    i��&�&	��0`��$I1dh&�~��=�4�OH4�G�!�!$��� D� L:�yб$��� ��`.O��(��hJ�!5�Y,ۃ�`�(��`�J�0\�I������ѿz�ʲ�P%J@
H  )(��  ��v�ھ�E\��8�`�[m��`Eq�
��Nq��/'NySJl�G0��E!�r�'
�$K
�����"���2�J�em��e��}c��f��1Ăi�����_zX�@��iMs@���#Q�������~�`��%I2S�%i$���$�w�I)$�+H����V�!$�I$̓9��'&��!	�}���=@��i�2����7�7��Cj����m�j�G;J_"8e�����k�Φg��@qۜ��vޓv�6�ޒI$q���������a�,6ʼE�Z�73�X�j���J��Jf"������l�҉7��8�ZPx�9���$�L��?qo�w�@��а�Lf%iuO;R4�7f�i����Z��[�6�v`�*q�oXx�k�I$��}�N{u3�߿f,v��tq(�� �"{�4(��¬�d�I$�Y������/S�]0ٸt52��^ZyU;N�����=1�]7MQd�I'��aޛ�̺g;QZ�n��)nѱ.g)s2�60ƕx�tXp_i�I$�2*�e�Bn���sn���.r�-����K"ZA,If�P�F:l�dli�m}ג���Qn{���.�P6HfدZ��͙�Lv�b"�ûB�.�,m�`�7K�J���MTR�p��Y�"�F33Z��!�K��"�F�����g�(4�{�{���`�o��lL!߹�\�4�P�R�ߎvm:�Eh��C�r2��Lq����`��L`����t��UTS%1DB�@ji(M#V^��2ց���d@���M��cё���c��ŵՓ-F�N*xזz|���F$}�/��Ϣ���6�V<��R�.�{@g��Zhs<�5!rU�K�m���=ǝ�+�C��B�*��Y,�5�T��S����+�0�/�C��ᨠB�p�hXs��`�mBХW��AĶ�|�
C�|�����~�x1��*=%Қ���z���/�,	�A0��)D�*]�by!��-�?\F�e�DLH`4�l+��*�J��]kY�35
BeE2;L��]�j�Sb�b�h�)B�16�E�V�!W�rEl7�V��*�+(XM���;'��B�����y�;���+%�21SbBZB�=B`M�;	�k9��ިhHb��X��
3�VY�	 ��mաZ�'
�}�
����~�Y8��j���jdf�� \I
%`��9�	��n��$.F�z���z�*>&%��� �v�8���A�f��0h��f�r�ZX		��cM5�o�N�����B�?�o*�G#"�xT.Hꪄ�C%V6Ɨ*k��qG E _A�"���x�B�����"���)�h�HZ�֗N��d�	��2�{�VlL��.V���w3RD}#�v�_�mh��.<�;FX�g���"�(H+�� 