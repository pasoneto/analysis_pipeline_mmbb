BZh91AY&SYz�^� A_�Py���g߰����`	z�=�͍z  ���@� ɤI15S���MO%=&���ɦ���$)4�     � "��F ��#&�!�� �� А� z� 4  9�&& &#4���d�#IF�&iI��O$�i�� z�4�5ހ�
�R�&�d�!�(Ao	��e���d��B
C�}YI'�z��As�����0<�Uh'ؘՠh� � $�� aL�  q��$�IӻT�WWkt�[���&5��$��<u�yK���f�k
l�%�������imD��Cj��ً+�1�-*[�>e���h�:d)V��U�3u���*���#��'uN��o����D36=jl���vy������kö�b�r�r�pGs\! )��ȠIq8z��ǻCh���Z��!��Z�V���J�W�U*��XStR$-ۃ~�̈́!10�}��i���B9YW�h�a��C" �1�2���[A6�dG�Z����hg��;;�3��#�t.g��.f�>���CQ��X��E�^3��'���2 ؝h�6U@��]�+%E����27a�p�`�DKv�GN3�dN"���m8ˬX�/Ԗ(M��n�ڝ��Ӿ����Gk[[w݃�#p[@�1��lc�vzb��q<wn&��N*�V��m�쇊<.��ӣ�}���Z W�ܬ�kLl�Ug� ��.ZC5F��V�i�č�WGD��r�4o*A��LY�F����U&�&��E�H�Fᨒ)��n��n71�=ք�=6�r��bv,9���&*����\&vŚ�6��:��1!��z��|�e##��i��KG���l&�tkVm��9K�3p�3*�0&�h���mAӝ
��Z�#��"u�-�WRt69i���Gh�%�e[_5�>�fn!�1+Je|��N�B涎Pf��W�C�-�pfq!CNv$�!��Fk	iه
cv���9���F�.��`��n��Y@x�Y�q`33l��m���^�;�V("#���		EN�S�G����*��G=y:h,�����7D�G�-A��D!M9�Iwd�$i(.ڐ.Ҡ%Ҕ2�B��ť� aG�n`��Ad��xk��գ�j���{�;�����d�vt[��	���To��Q��U�C�n�����n;�����wo.;��K���&G�w�w'v�q� ��b ?�R4�5?���}�BrG�[��1��㦞��-�qTMC�b��Н'�*���2�SI��$��4��fy�P�̡��q�V:Q�^M�o����/��lߪ��o�" ��.� �G�Q6݁�9w�׾�D؞��1�j��� ��1�f����qwt�s���RHD�������:!a�M$"xvzK�Al7��I�R�:��bS�3�A1�|�aS �p\�b�3��6��9��N����f�f	�7�Ӆ��̺�H"��i��:���.��ˑȭa��\�6���;���6w]ϴoDF��e^/���\��`2/[�3jx5z8��Mil���+2ɕ��l �x2�[����h�%ql"=�p��a�k�Jǐ{Nc0��:�҄�ӫ���6&��ŷ�p}4��/��ɽ��9�Ґ"y�'��/�!"PPPX# �E�������EA`�A� BD�xv�5D�7�0Lӓbɯ!0dѨ��HaW,	�8�:�,��~� ���c�J5�G�I���@DDqw��Y��������`R6Pp��zrss\�Cy`�d`���6V�*30��Ui.��E[�.r"O`�py�A�E��쑩0/�`%)�{��"�(H=E/M 