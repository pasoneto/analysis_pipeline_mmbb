BZh91AY&SY7J< �_�Py���g߰����`
������1T� �����k_t�I"b �(�z���?Q=#@h4d�*z�"B&h �6�` 0"��ꪛS@ 4hh     ~��h4 i��  d  Q*y4F�  4  �DȊ=F���M�3Q� �h��iR��0 !(��� ��来I�������jL�_�ؤF�4}lqrU׽�$�R��D�TZ��ڹ1�S#OW[*/�n� ��R�P 	(j���R@��ID]�dZ�06DW��R�h�^��X���m���������R4^��iW�x ���O��W�z|H�ɧ�7;�4Γ�N� �K,�p��V?s�1���< ��Q��B�����eC��jU�ƫ�~E*�Ly���&�R���C����%4>��y-�Nn����.{oO�<�1�@���d��e6Vr���UW�9�U]�>h�g* ��e���3&"*rgeL��	6��Ɉ���UUf]�f��Ȉ|ʝ����xx�4��a��M�pe��g��U�RV��xa{e,&l�����)�E*I҄�C�j�O�Mz=�z�E��a�yRE��" �H6A�͇F��GG�h�p�]�����Ҳa�{��Mg��Ť$$�B֋�0�.��������eNڡ�ַ+����[U�6��8m���r�L(ҧ*�4m��G
`�{�F����!�w�ޥ�+�����Y��d���VoWw�J:x[��QjwS.9p�`�B��GB6"DX�
[��Գjt��2�ö��Ka��v�6�-�^y����uT�UU<-o1ᄝh�I�$�I�<Q#bZ�9S3���M�vvvx_�N�sz�.u1]���^a��w-�3���8������$˦陶�G�IZ�΋(���8�i��"K �0��(�f(�Qn"M��k����3�TTYئ=av��E�H�t	�r��$�dX��8�� ����F�wk�C󛈪j������BBP��5A�ކl8Y�F6O\ p���#eM�:I�8B(c(�
89���f��lB��m^c���P���Ĉ�R9$�6a�"�)G8nr��m�Xw[�ktwp��1�[j"<���?d��:(�vI�\��a���J�$�E(�e��{�Iދ��r�0C���}Nfٷ��{5¬�KIX��l��lX8�l��,�GAg	<�0F��i����U)JR�{iUT�H���x|��ܛ��q���2�V�a�1��lhU�--ib�����E�%*Rb��(QrReF0.IkKX��3Rc4�Lc	�U/�5
S�2��S���/�H�U`�[&�gT7O���<	�m<��j�|���No~�*�\�A��-���d�/}���au�`O�����P�c��o7���D��B�N{�4)�%9`�_�r8\�K1��IV���z��k��� ��àB� @��"@���9g3�RLs;�-i����ꖷ��O���
��{��<����
��o&�Y�ɞ_�8O��H�c��VZNZ�ê(8���J�,��(FV1hPo'γmt�۲��,@�B%J
�U��HO�n4�_��H���'�.�wy��)��x{��$%?��-M���)0��|kV�{�jo�L2 ���p%,X���$a�As%2P
�QaO��G����v`h������d(��$���9�0�m3CǏet8Ԩ���������a@��RX�
N�ٍ�بh�HC�c�.d��;�'t�Oj�t������kiej$ËC����c���P&@�N_��VH:�#�N�[�|��Z��"���4�Y:g�6��d��)�R���S�}[      !               	  �+fnL9,ʩ*̪��2i:�[)��T���ꘆ�1R�O�õ��W�#���P�dQ��XNPBBP\d%^��D�Ҟ���]���y�x*Zp�.z&�˕9���T�pvpK�}�����s	��x��d\�@��˾�25)��9��0$�[�a�.�p� n�x