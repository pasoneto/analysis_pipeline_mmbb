BZh91AY&SY�4� {߀@y���g߰����`	9��ϟ`%�U^m��)�����F��@� dh  �i� 20  14�T��UQa24`A�2h�d����) �&�CC	��  �AFS�M53DچA���4���dj���?ToAG��4 2=M���W���*Q��Hh��]A����v�#��
�@����*�D$�B�o��g�'��@H� ����$�  �D���J��#u�ubyP��%�󹱙�'�[AX�"��Zhm�bm�A`�`(.2s�����X,-q>'�����B.E7��buɌ��Z�Uj��|�Tk��9�s3LӼ�:#��D"ES���T�����r�p�{B��g����xZ�	�fz]!ʏ0�Wݛ�Æ�o�=d�&tѭMU0&i��@2�@	� U�U�@ Υi�
T �ۺz��ؐG7ޛ9_d�&hw�,!�f�\ڑ<�����U���&�Ax��D�L�0�1��\���f��:]]��(����J+���hZ`mm�,��,����˙k����SW��������,����� dL6h4Pli�V����KgN[0v�X��B���"����m��ךᰒ�+4lW�n�L��$U*�,�N�Ku/l81G-��q��l�iV8Z3�$�w��k85�^@���70 �.�ҫ�>�� f�g����5}ZR-�k�`��K%� ���I�8�7�PL6Hi0
P����<Qu�,:�F���@,9ۀpp�Շ��[���& 7�e�g�zZE�U�[�Xt�MK�9�c D��jJ(2��N���%� �XDf�BW�08��R"f�@���� 80U��EX[u_af�` !�/O��&Zl	
t"@�t.���� Q���h
\m�$r�����B��-{@8%��g�����-k�,+"��	��q�0�2�sca�,5�(gA�ƃh�@��%�qZ�c�<��K�5�8��?9�6��1�sm�4	(E��_��\�K��{,B�VR�- �,�!Z0J �5iJ���i(�GkX��H� �S�&�b�Lf�\�!����}���@��N��r'�R6+�#
�� ߯6��~'Om�~�A���Kn��=6��
(,�5iKH�B,�89F`���303 *o��E��{>���:4{����r��ۡ�A�4b��hH����}*��8��Q/�ēߤ������rlb�]�i}|2����܈T8��w�{�ʰ�3�#P3�{��^�ɫ	 �!c
,3�@I��Q7�a����9q�h�o'f��*��E�a�%�n��D��i�%�z �a�(�2�A���p�t�.����sJ�A
�3�X�x���_koa���ڰ�QL����0 ��
Cx�/�����3TY���X���V����(P%E�s������YMu�4>�C@�������cSL�o�Q� 4m����Y3BG��Q��i�#����r!#�}{F(f�!,:B�+5�#n'W�0b%�UQ}�B�:��Q�
��>�������OW�`�
���60n�))#�r�t��!Q�Y�-�1�VW:�i}0`����!�0`����$�ch`������;
��!
$L��V��T���XD4Sf�Kd��H�L(1�b�H1i�T"��(!�����$��w�N�A���5q��u(^y4h0z���� �"���U�����z+<�0q�D_b�h쭏�G��6�0��-?��H�
�F� 