BZh91AY&SY(>� �_�Py����߰����`_��e� �+���0�)����=@      '�RT��P @  S��USA�4b� �i� � FR�6���  0&&�	�&L�&	�����F���&���~��4�j yOL��y$O�jH-�B������L�+���Ns�PeR"%K(��<*��р�g)�#�E�FU4ׯ�zym�6�A �	@J�$J���I	@�$�Z��`�:�`�d���?������l?�\�'�;yK8!�
�C�k;�4��jj|�Af
|K\�NbX�-\�LdA�`�:}���>4��B��,X�ZV�k�ờ�nױ�u/x���j�	����o��n��:�7n�x'H"I$I%��2�%0I�$���$�I:I%)%�Ϋ<��Nx�'����D�IJ��ï���ު�ʍ��/�C�/�ڡ���$�L��s�gz^,�h�,�N�/L��-br�L�ݹ���#:�w������l�� 2�LSz�$C(����C(��Y<�<P1w�/�&�b2�ژs�	W��aA�3e^@�&9"��o��[�9v{Gb(��m��%�/j�Pl�l��"�Ⱦf������h�[V�w�Pn��{�R����p �R��v�U�Z�$�A���\LJ�)�So��*]��*ɓ9'�q�bf�^h�̲I$�h��Y�Tt�^�(�]�9[	f�r���$vdr�a+���m�UaD�I$7�U���+]�!�v�J�����ʉɔ"{���o`���k`��I$�cZ#!	��(���r�-��W"q�)\;���ڨ�I�F��O/��V�� "���&!��ޖ��d��U��D  Gx������8cWV��&ҶL���d�:ܖ�6�]   �ɷy�]�j���v�`���d�͍Ŏ��%HEW����%��^��Y4x������>�F1bI���
*� @�ޘ����ZQR�*Z��劔T��(��)R/z�W�Z����0&�d1�ȑ2%L��	��Vja���TƏ[_J�B�"U$�M�󰎏��L+k��r�r�k�����㡜��,���q�$�+c7I�uL@�w��<���/3L^���D�?�����[?q��L�ޤD��R��F��X{�n�z1O(��a����T�C7ˇOz"}�&�i��ZxuY(w�$��c������3�`�9��"D�uK�c{�C��*�yd�P��v��RC������{o�s,ƥ�v.��]K�>��Z6��<['3"E��(T��8�l�4FOZ�O�nSs>�j�7%,���nz��W����±��o�JDK��6��s����YǬ�O.��F�bt��u���a��y���mu&�S�GgJ"]������<�\�b莤�8�$�Q�=���������4�,�4N�W���.t��u��L	$��e��?{��3�X�E!��p�1z�X��ˆ`�v��Q�k*2>)"Z0g{���oIUn(��;��T����lhO��pl�#����*�m��zex'C�ĳ��0��jM,	���*Tu8�](�Μ�~3d��&Q�w��Zኪh�jz7KI���+T��+:�G��̚W4j:�Zr�����u��_��47M�f*�VY���ѵRɋe��t�����)N�Z�ȴ=�	��m�Ԕ��=rO��9ٺ�)��M�ӎ5F��Ɨ��ޤ�,to���)�@��