BZh91AY&SYBM�� 	߀Pyc����߰����`�8ܯ���
( � Ѫ(%�cNz���iOSC&� �4  O!R�A  �  4 �����=   =      ��U@h  F�   QFD�� �L�z���6�PL��SH��JjS=Pj#j=F�� �3� ��*
 �UP/�y��j�>[�	O�̅K����'��%���� �
�%$��I}I��.e]\�Ue� � �*�@( ��  UU�z䗒�R�S!k.����$�Ơ��]y8�%P����E�n�zJq7�8�ț�+˽��X4I�64����FpB��*��� �t#��5p�@��������T�&�I�^�6es����{���n�C7A`���0���-911�.�^����[$yv�|zt��2�Z:l5���V�P3����ٷ��s�>N=�9ε��\��嶜ECl:m���i��!��x��x��m��m��6�wl�	6ӡ�ź7�����9��"�ӑG:�� YWN�!�}���4#r�L'�ε��h�Y" �����$��j���K���Əϳ�����H�f����L��%���n�2�c��8����(���
U�*J�oӘ�L�f��X���wrYYJR����FeXil"���Ĭ�����S�R�$e�M�G�8�x�\���m�[Hex��e#�>W>��s�<�6�(���sP�E$���07$�L�;q�"!�0�Da|jN������!�i�m�[,�A�)�GN�d����׀� �h�����1�4b&�r6��I$��ӷ�tӧ���ۉ*4��6��\x�m�ێ#.�In����M4�n�v׵+�1�z�]t뮺�z{��wwwws��4�m6�-���N�zC�4���n2�m4��-�e�u&�r\����4��,#K]{�����X�n�onw���������(�Zq�2�o�-6�(�m�2m�m6����ܜGå��ǌy�<����m�9�o�/��'�x������'��x��4���:e���C�m�M�㥢ݜe��!�pֵ�iTȢ5�R)�vF��N:i��ݹ]�]�#�;z��xx�6��t�������{걢��H<�$��"����vD��6��YvÝ���fM�;�N�a�[��Gim/kt�v��q��ws��I=ZeoN:Fޞ��N���'�]����\H���6�\���~�ĝ<x��t�UߒG�����r��}*B"%I�Ą�U*�_���G�co�-�b���[̮���clEt��\U�k,JA��t�JJ0��!.ňEB�P��T!KY-YE�Y�V-Y��c��.*Ն0aX��%f*��J�i�$H
���F,
$B��.hH7Qi)���΋���v�{��`	D��Q�|��3�K��x4���k��y&P��q���=��q.͆�{:����58$ �0�{�&�ܔ�3�KpL�; �� �2p�������+��&���J���-��� �A�;�n;PG�m7oT���I>��|�_����$�]J��Y��^�K/�~��c1�]vL.؇Apk��k-5�ѶR���G��/�Q���!U��v+!J�貤�%��]�!Q^��_ewGG�������@C D�]�90T4ȷ��hu��K��Pv��g/���P����$ʨ1���m�xR��BF����,��y���wR�c��V܂@�E��l�Ŕx�ƅ�Pc3�r|�J�`���Ț�*�������7	�c ���zOh0�#�?"���!�uU��~|�*��}*��4u3U���Aa\���+��� �F�5W�4�W?����ٲ�^�\J��[�r��V���Ҋ�Q-���׬"v;PG� r��� �a��>��(��@3���6���p�6<R���_C'��qY*���T>���̛��d        �                ��jK�?���J���)V/#bU�'h�ģ+0�Z�A��Z��nl��0����!}�vå����j!hp��/�nu.��R�&f&C]���i���0?+��M5_�#�x�UJ�p�!oq�u@�'&`��t9r�2�7�-� ��1iw��y�W�`�ID��"�(H!&�� 