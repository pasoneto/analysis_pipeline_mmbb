BZh91AY&SY��*T /_�@y���g߰����`	?z�{��s�� �\�  D��T�M4zS�2d��4�Ha`�&�"       *������     $ԑ�)���4�z�� 9�&L�0�&&��!�0# � A< �'�Ojjy�A�j����4�����(���D�-XD���FX��PHD3C��%W�2E#�@&AO�H������q�=v��M!� I�	 ֤�  �H$ �� 	 I��kZ�{���8�6�>���s�kײ�E�J~��8
�mAP�Cm��D�Q*��Z�������"�n�	Fx&���F���)&g㷍ZչdLE]ܻ����Ϊ�9wUU��U��,����hA��bI���<��zu�*�����\	4��-��՞�UR�V�*�걌�j��1�/u���bꪷ�j��_,R���\�7�v�y�	�"=�l��>�"0��28��YP���� �3α���0/��`����Ũ�B�t��l�-R=��R��D�8*u6�c>�{j��%�2H����ċ$��Q3���A��8����bڐ�UV#���8�#)(K�C�LU`��h͋*���2��+Z5�m�H$+0����l���3��סxbX�a|iJ;`+Aؽl@�[l��I�+Վ�;��k���v��P�'�D;�qP��9j�!h�/��r�-oj��h^Gt��%B�Zd��]z�Z�+�9��!�V ���/e���9��\cͲ��UNƮ��"�/}v�H��LLdS�$��ؘ`�h���2
�H+V\Y�k�\8@p 4'��J"Sm�V�ͨ+�^��ҕpx�9�h^.�mƢ���x��"D!��f;!��� ��Dn.��Kս��+�	���c�J��?�`P�
WcxI��4u-a���l�w5�J�7a���u��=�=f�*�.���[B��ɺſ'���I�!��I�@�A�UU�BQSŜ��=�%�)����Ie�(�аbO8E�PdD$��V�E(&%�(�&%�(
��Lք�e "k��^Q*D3fͫь E��$M�V�������lr�,�%�ڿ���)�~�� ��4.����.�е@K�m+e�({�8�i�I����HK�(���>�/$���>��3{�AS���������^��!�2��p�~�h��._ Q�-y��!Ҳqı�?�� �Y-r�He���3�ĠQ��1���!�0#�%��S��['���KeT;	�*HC�7R��	r���¦Cb|��c`��FX� `y�f������>*nt����0���!.wq�	�?N�� ��	! �G�J\��������.����(|��Pvh=a�,���a���w��M�(���1t���Z�Ð�aEx��C�S�v�����\�`�@��͝�gu7���bA׺�a������X�$��50 ���!�@Ndd���`�F�@*I����~�@Ͱ(�B�w�Gy�P� X���m3ǽ��$��>cb73�� ��"���Pݨ5d�Q�5;�����,X�c ��TAEF ��Ł!�a���4P�!���4�lX5�K�P��(^h��si<����=�eAƃٹ����·״.
8w���Z �/&�M��`%Cq@=8rr�A��hd\#�l-�#ho�!�P��U�duJ\ә�H|���[���[
w0��?���)���R�