BZh91AY&SYvE�� �߀`yc���g߰����`?���:���v  (��zjz�P��4 bh�	��? OQT��2 h���@ M?�UI�4b2d��C�A���00�!2��A��   �& �4d40	�10T����4ɤcF�6�F������z���%u�.B#$��|^W���	3��_.s�[���T	�T|����Ō�&�RL�
�T3�����>���Ǯ  �   ���    GD �.��Xp�܏��Ѐ��u�GI���(�d�J �B	1DV3�D͉��O��!3��d�(7�j#A]�eul.jڜ��IXq�
s� ��	�=�b8�	�A�((���9��97�c��A��i�R#l��]gb�|~f�>�~mz��A����USom�m�m���a�i��m�n"!��a����p�f.P�x�}�:�t@ {<���@w��& �	�f��`F��I ����T���.U� ��$�T	��׹z��z�dQ�M=p65ț�.��/u<}�Ԑu$^־'u�"i��m�� JJ��I#!����q�H��^��ށ��T��V+)�eY5 �f�@d;; ��[�
�d��c��m��v��H#l��,фN���6C`��_�(a�J�����L�e�9�ZZ�˄�fҸt����E���I$0�B��w9őWX9q��;\g`�y�1� Ь,��G��m�9)�gp&�]\�v�e��c���kG2�ֳ`7���܉�I$�R�tvn뭝Vʨ���Z���.pT�)��	}O24 iԊ�
šæ�I$���+�6��ӫ�0Z�3)m�Q��$n��%\�ԓ�c[w"�bt�I"PQ�b��6+|�����x��WɨCT�Ge�I&F��� 3q��щ�r"�E
!޵�X����E��I&��Sp�F�n��dA����8f+'[�8x1�	A����)$K\����4��d��|��m�kV�0�d��)�E�(��l���QEVt��K(¬���*(��J*I�ケV8R\�a�������(���h�Ls��Mjc,B4�|+�)		 R'wA���wf0ب:�:W}����X�������̖��%"m�*y_���ߢ�86=)ާ��w�M���n��'d��=O�{���2�7��k�D��e��ښrϹO����$�Jcol��������̑>��i�6�����N,^���ΩQk��=��k|��:2\Lev��^�9��sS�u,����S��	���z2�*a|ʜ����[O�n�o+'$~����l̑r�T�R���OC�i��������UM����~���>�.��.h����u��̿9���ǡ��RTi��4�q�Væp2�3#��5�'f\$��Y�TVgվd���8ƹ�s�"w=)C
�;XTݔjVɛ��I�a<��&�'ѿm�H�P��`�����!lS6F�%�k���gݡ�e�S�F�K��� ���U���g9*���H�y�y���-I�<�v����-9x�{q8��[庚Jw'��[�y�3v���$M�`�:�J�N�{��5&�6���:X�Z�E(�H��&�N2��%4�/��jȉ�T�՟#F9�gC����G3s�*��wnf{���KN,�8�N���ٺ�N͌�p�1����o�����z�.Y��q�g�й��ʕ���O�[��X�RT�������H�
ȷ4�