BZh91AY&SY
`$q |_�@y���g߰����`�����d�2 5@IB4Ќ��B�z���4M���ҕ45`�h`h )����d���40M0h�0�Ȁ��e��=� � 9�&L�0�&&��!�0# T�4A1��&�4� �di�4�V	"x�AH�c 2���q`�%�)�#��G����P-�Σ��5Ug��i�$�P�j,�eSE<�=]�X�� ! @     D{V�t�ǍI�t~G�c"3���(�<��G'Cغxxl��^�m��a9w ��)��D(.S=؇,LP&hu�q5Q���q���:�������$瑖�]CY��<�_�r���Li�8�y����
oY��A$���2N�I$�I�;�I$�I$�$���	$�XʒN�N��\�����J(�y=�����U`z�l�zl�[�m���"�wl�P��$�Nr�YQ,�ʫ�Ʀ��j���/�ص|n���6���"�sX�4o��CТ�卦�h/u} �Qk��(l,�������(��
D�u���p��J�fpS#�Y�@��y�K-�T�D�Q��<��Ka�y��i��}M�T�ejÃm�~�e�(�W���	U�̌%Z�J	�ը���X�W�vm��c��՛��S�)�]�ʹ3yP[1��~%]i��H#g��Y�I��m��Q��oh�k�|����%�)�q��.sa���W!=�GaQXI$�k�l�x�.��c�jm�;W ZZY�.gD�i����E�	I�;O�
x�P���WL3;����|��jWE��� j��k4�69i|�C6�|N����=�O͘WӺ  @�w6�h���a�E�)r��52xw�3q1�k�\L  Ϗ�BM���R�b�ڐSs��٭���Ύ��k�=��%B�zI"A1Ǟ�|x0ǚb\����r�1IrI��d0DQQE
�IEEeV*(��R,QEQEQEUK+`��4�dL�L�r��1$��)� �*�	�L
,�~��%&įj`�˛���A��ID��@�������ў�X�|W���gَ��O��Ԅ�tͳV�؊4��R�Z0�3�/��!dO;K�,�-����-/�����Й��zZ��Պq��	���S�=�<o�>Q�[��M��ӻ���G��6HD1�aL�|�C����a�&�c�=��٘������-��������RC�Q%L-�ZT��,�f~͌��l�#��5�y-*!R�J
��}&Qwyn��97ʩ��o��4&E��s�~��yͷ���\�v��K�3??J�s��,dq����:�3�y��9#O�yo����4�����7K���#��8TD�!�z���w0w����Z�M�
M����R��n�c$IC_n	��Ӿa=�B�)�j��X�/6�\_B�z�,�FG��H��Vv�z=[�Un0��0Obj�R|�c����v�-4�M���W`Ǎ�8�A0���Rg2���I"SH�*t8��<"r����{+�^g�Գ �PH�BjOk����c�[L*S�n�ӄh�tih�{cB��Ά9�t̡7+se�*ֳ���ѵR�uM���ɛ2��S�sJ�>ldc�l�i)�T���bݡ�ѓW���Q�1�ݡءؤ�5���ܑN$�	@