BZh91AY&SY�'cd �_�Py���g߰����`?���Q�H  /
�
��BI �jz������@ 2S�i�jm�D�&bd`��4z ɠUO��UT �#M444��h2h41F��D�� Ѡ    sbh0�2d��`�i���!�D�hB�����&�O@���&�h2���ie��ȈR
%�@��4=Ņ�0��;�u�� �B�`H|0�|�WS1H���(��9ë���Ën���9� H%4�LM �4 �"i I4 �Z��j����(ׂ�!$3Dzccg6It�sGn�:ynuc�����ʵ7"K�C33
{�2��8aOC����*g�f�
R�hB/hQ�c��[�u�5�J%�ZY��JIc�7�Ϛ����j�&��;
�,a
�82ς8�V�1����5*�ZK�[V6����b79Ұ��[l�6��8�� P������9�Ǌ��O��ԗ���I(��$����IZ����|���ZX�mwwb�r��IUZ�v�7wmU3�5��>_�����a�~���o{3é��h:Y��h�T j�>S�1^�eg,8���ĉh��Q�jV{�
���Z&5K<<<��!٢���+�b���J���}󃝁��JD��!���|�̓33k��JŨI`�M�%��E!��P���LPa����,����r�2��&[�0J:޶ccq���XSTβ��J[lQ6���Vi20��.|��^`9κ�ޣT�>x�ȇn$���m�	$�H�C�sۈ�%���۾�e�{�F�`�"y�(�)��6�N��ikF��I�7`��h����i�V#Dq7b��Zm���TJp�fn`������;�-�T�Fwɫ�I$�Ȑ���^Fؗ\����°�S��O`�/��ۡ��Cȑ9�P�����".�_)�L4��a�*�T���MGZ/�ӒI$���bf���uf޳��l ��S������}� �zr���M��a��2��<Kc���v��4q^�����Jx����6�$�I�E%߀�OE�`���ǐ^,N8R���0�
Vѕo"ҝ�����ga޶�,���Υ���8��I$S�B��	�-��gCc�l.^'x�.��;��1V�B�+��R�0����E��.S���7�i�[4�+�$A$:�׏;b-㑔&���k,a�u_*�t2���k�W�j��y�/��I�ym�C���0%�8��p�E^H�����nn���(�2P�4���ZFא[(Z+f���V6$��k:K!mˤ>�\�}�np�ҕ�b�����T�T�
�^�s5�����S��kC3-�:VcǢ��X�����a��	��͝�A�7ńDE�E� �S�X�R���r�g��QсE�6-�#q� �$C�A@D� ���HŪR�X`D D A��A��P�fSc ��I�������R$�!�
"���8$!��%-�Y׸��"2	3%{-�q���c�IJO|�
q��@��������)9[*���/O֥���q#w[�(4��zG���4<ǜ�o!��x�Gx�{�Fӗ�;vz��ٺ�,G�� P�[���1D��^�7)��F2H>zl:D���I*��h�&��#1��r&��-:��ٮQ�3�rܠ�s�e�^W9yC�4��cC�g��W�뽇�|�A[X�NE)�@�$h�F~��ƙ �	���[���P$	B0� V�,�G��hW1�S�ը�;�F�����Ci�
5��<�>B�3o��( ���(2(���o��9w��	�Ҵ�8�U��A���B+�(%��,�\��Z�D��Xgf�c�;��Hn2q�|@lyb*�Y�� �9΄��Z<wLɭ��HYޝw.q��m�ĸ���Ïϻ��4|K����aS�V �ٰv�#�@�Qʨ���n���HX����ܬ��xEG�,��:� �è��z�R�8k���D*SaD�P��-Ã�ǰsL �jo����tQUUUaUUUTUEUUUUQUE�QTQUUaE��QUQE�TaU�EVHB:Ap��0a������`+�Fe4�'=�ը{�b<�h�>W��D�x���RbQZ���!$*K�Gmɘ�P�L�������S���dff�9�
���k.&�	��&"��|� ���>%5��"AvF��~�,24�K��Øe) �sّ���"�(HT��� 