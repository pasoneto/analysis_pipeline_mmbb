BZh91AY&SY�3e� k_�@y���g߰����`���( <��C@ H�M4D�mF��L0 	��D�JE  4� h  �~��i��# �CF�@��2�f�=M��Ѩ�4 Ѧ�9�&L�0�&&��!�0# T�4�R`���?@��P��`��yOS�f"v�
���y�'S�/Lw?�2-�*���)���_��͌���I2T>��*TΞ=��7�{�߀� "�(PA �	   D$����t;�u�9c��Fk-�%�5��i�=�����^i��R��!'q#"�Pƞ#!���]�Sj���8�0I����OwX�mA��F��Qm�]3�І�Gm�y�dЃ��@)��H"�H0�XJ�alO�	"JI:H$��K$�)$�IBI)H$�ID$��I'I'wt�&�o���}��u�ß����5�`���~�x_8�W;xt�u�m��՘��V��7��Jy�F8�o:�*�d�O]&������3��y���rI�7��W�Zl&�k��cuy��F�Y�&�e�ҫT�OG���E������9o��ƚq�`�ô�I'*�(�ݣ��/"8T���W|Koj��j-0��
�����19Y3ԇ��hgt�}���[ȑ^ō-��$�Kgl�g���l���Ռ���o����V�ˉn�$�]���L6���L�dK�$�ILh;O2�q+@�9f�KD5�f�Kd�D+�z@����(3�kD�I$�����.�y�m��b�S�Mmb�끧)���5+��h�XI$�L�ٙi};[�SH�`M{��ʷ�)�6��]TSn���	���@cr�ND��:-����b��u5tǬgZ���&�4� ����?Xbi������M��yS@ �EB���%6���ڷu���km:�o���M��5׸>c�6��1���bb���j�B8�<�!FJ+	x���J*(���(���T��X��(��QEjF+Q���E��1EUA@�D EC 4,�׈�����D5v��}$@�����ɹ�?߲Vt���cq^��g~x�$Q����l��{Z�a�EG��n��Ξ���=�}������ɽ�"s��ὧ����,5L��"�hY>�նzT���Ўۦ��B��t�|T��M9��䎁��gqr0��?~RǞ;�1�(E�-/F��=�u9܈T8�ck��C*��ʥ����}��>u1b�'�Q
�[�ZT�k�Y��^[�9��d���mȐ��R�J%[cWY�]�-�y��J���r��3L�x��e���)��b�O.F Y!�k�Y�݅	BJ^%*a!��2�M�dм�LK��F���&�A�MQY'u_3H��M(�4=��(r�zVz�T�x�[fNF
N��u�%�0��"Jy��|��SY���L�)M�U{Ռ2��6��T�(��3Z�irD��������ȕV��"{L��6K)>g���~�-5�M�xybiԬ��0v3����u�Y���50DJf?��S���='���keez�S8�ּ�.���v��I{a+d�an�:�N���ׄg����.��k���un���-��ڭk72��8*Y.��,��55x*�+�ׅ��c#��p��{$s�8jih�_&�O�%�Q�1���ޡޤ����EܑN$;�}@