BZh91AY&SY���b <_�Py���g߰����`	���Os�r  Y80

d"�!�2�e��'�� 4S�h	@��$ & 4`L# ��U 4 2  hd   �QM ���hh=A�@   �4d���`F�b0L�`� �"a5=F���D�����i�W8��t�!!DK�P<�9!�B%�}�K?c!��풫��#�@&L�H�����0��w�4�M4ﺶ�J�n˻��*�T T @ Q  ,��۴���,�ӱ�|ڹ��uq4�u��mf�N��p,�DJZ�q�f�>�3���[]7�N&�a�ŏ�>TC�k�S��oX�w9cGQ�������Ϭ�w���֢��-:�V(Â�V�����=s�u���7=wu��#q/��Ӟ����ZK��%�'B�I�UU�VXL1��l-�-�J˃#�
�F���F���h����'�Q����N��H��'�Rij��x���9[TAi#i��h�Zg
�;A�L@��N��l�-�G�l��M��0�&BQ�3s�S$9��C<�M�M��=8��_ `�5��$�嬁�����;��N�����D��U�e;�������
�-`V+��W��ֻZW#��%lQ�M��h�f/h����u�<E@O����6{n���Lǧ8Y,5�˱����]�5 �N��c���-�B'�xn���r��f�-�N[[�r�	YJ��B64��(A8q���� ��513Y�Uf�ep�0-l+%�
��v(��nU�ҽb!7&�EY�%�+��WhIšh�W��D��Nx%NБ���ؼU�Yy�'o��)\���e"x�e���Я2�poM�;��8рgB�`�Bd7DTO��А@^����s{�65FRͨ@�BS�Д`���G@/C�����:\h˦�f	z�s���	���gݛ�7�-�/NGA������UT���x�p�Jdv��i4��I�RYb��4���|���Q�.`��D�HK�#w!tʤ���
v�BX��2��%H����b@��""!#��V���)���Q�[��^��?�a���d�~s�%�@ɪ��1�ϥ�<u�iyv���|��!I�;N�D��R�Y�7�&dQ��ሺ�jm��w�HT�a � "�����3��!�)�2�whD�[�D~K��D�u�������m ��Y�r�8e���3��@�1�e�ze�yHݺ]� %1�y���ځ�TW0�z�P	
O:���'5.@I`��r�S!D֟�1�i��a@��W0(�	����w����N0�AD ��	�k=���S����_rHB����4^���+}���8q,��=sX/��ֆ��|�y�3�ᱴi�|W�**#Ci�� c$���r����@��8(���
s�Q���)�˙��F �
 �gh@��M��UlH:��M_8T?��P0�@A�1�f��Ϣ�j`���̡�[�x�d	���m ����e�������PȐ<��fo���H<]}�#b9���` �{�"��z¡�Pj*0� A��n�rH�0X#��c ,d+ Ȋ2,�"Ȝ�*L
$7�̓	�ذi�.�@<�P��`#@��xK�7s���C����V��<eo���Drv���Y��3/���	Bƹp�8p6y���������9�lz��9]�7J\Ӂ�$>�A	���|V�`�?��H�
��@