BZh91AY&SY�~� s߀@y���g߰����`���ݪ �\MP6���O5��Si� �� 4h ��@j%�M22i�@ O��UT�a4d`A�di����)�50@ё�@  4�12dф�14�&�JL��b�i��2L�i��A����i�e�����@� �P�?cyp���}!x|���
 �0�����qPE��o"��"�yxs��.�Y	�� d��   �3�X��Ȫo�>n���T�FyZ������@�`dZ���u��!CõHw�^ٔ���=K10m�k4�i"�3,�!`��o	��-2�X�3-��k���6ђ_i���P�Ũ�	;^Q\���k��}h�,��Du��bE$I����)$�X�"JV�I%	$���I)`�R�$�$II%v;{u�A!<�:����Ipz� �R�6�.��$��V<)$��&m�pVWRqR�N��M����UyO ��� óZ�և$4im�X;�	Um��l��\�;�1:T&�ɓe�#" vx0A�F��f�{�
w�1T,0�\M*84R��1e���(����{����<h�[�9F�m��w�MB�h6U����+�4�����
,�A�:"�b#	$����E�b�Yڥ�CCT�����KHn���̧��8���[�-l���UZ�;qT��ũ�hii^��m�%��I$�]h�x�殟Rq��)��ź̺vm��ʉg�n�$�I,�Ju����ඛ���/x�"4�R`����*x܃"'�*ŵa$�$�����f�׻�#����6�8kC����Ev�{�g�2\�36��KU�0ǂ��g�n� ���Ba`��I�$���e-���ݾ333M�g�����v/�rwb��"��[�1����"7�)�Em�;��{���}�ѓ�R�7:���<a�L0���I�!�;�9����a�%����A�RX�na
 @�����
��J @��$Xr�!DCfBHM��I ��`�""���V�
$m��yD�BEd^N�6F���ϟH�#U�pWǟ�L���^s��N�����o�(&l�b#8�R)2��@���*1�'/��Bƞu��,�.�q��T�c!{�B��4��=F��s�w��
������ �g�~#�Md�a��/J=|�J���d�"�Q��.Hc:dpTpD���/|�à�F-���F����'��>�s0DD%� �F���Pe��	8�� ��®��J1�0S#zX�
t�C̎��nj0�o
y݇[��t`�ԠD�*f���<���w��0߂ľ�o��{�9�ag�*C4��|��d��ƃl�/���-]�i�2s����Ǥ`�9�\vGe�io7�as�{,X��٨*��<n�=[����,7FF�K�*@[��ip(�2$�ڂ���F�P%?o^�d�f����j�|�r��̣��ug��g�����p1a�9�R���j��8�Qh��y���r���|�C�'cg�1,���1=#SR��C �n�U%z�s�.C��b���nc����Š ��M�eh��f���`k#A���y��X�Hm,!D<
�_a��䧻�Sf&�%�Y��=���M�o�bt��S8���)����p