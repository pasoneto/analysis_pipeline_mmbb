BZh91AY&SY�� t_�@y���g߰����`����D���T��)B)SL$�)�F�����CA�i�h2M�5"��=@4bdd�dbh��S�?�T��@1 �����0��BSA�@44    4d���`F�b0L�`�$�	���S�yS������P ���OS�v
�
��?FI4�@�X,�G��	@$&�א�6��T��4����
5c�~���t�)JD� L� @L H��P 	�E-M+�u:�>C�Vc�-�&TÚ�ۆ׻�����o�td�'
r�@�eA�A�`�@�,�Y@�L71Ky������O�;=c��;3T-ķB�H�	�-H�K0�}i^b2�� RV頉{3`˓���[��^S6YU�"�"�%r�I%i�wwJӲp�KI�wwI$�t�J�d�;�K��v Q���W�2�DÖ�^�i�*�ycTD���f��66�LLLP0�ל���z؈8�̂����k����@֯��t���i_Y#mނ�[���1)��0�,�9�=�_1��:zZ��Vi�Z�[g%�ɬ=�U}b�W1�3�w�)!$�m�]*����})�%�'��'��+f���BGrF��0�h`S��EQ� Iz6il�0�2m/�ıSJæf���x��9����I,C�<��ꇽ��[��8�+1Ƞ�92p��hi@V�bhQP�I$�I1OBj��Z��,�d(�5�6����p�O1�g�-��I$��nn"�G4�����;��i�T��Ia+����"McmPI$�I�x0%v)�X�ˣ[GY���I�Յ6w��D�I$�jJ(M����8ܵI58Rk���w���Jr$��)�&
�rbK7٪�Ԫu`�x��e�W5HjgxH�%����!��Q�Ej]I�y��eK���ʮXa���o0�8�61�m��Đ�������aB�K��:��`�����L0aѐ0dڀi�N�L`�`�4Ɩ�@���%UAF\�(e���5�k�S�e�!��̿AI�l����}���+�����O���h�z��5}~���	�ǃN�_���$^�:1r1�t��X���2=���3!pU�N]�w����D��@�s�rj�b֙$E3N�!� ?mZ���H^h������d
�$�ϕ�[�,�+��BcMN�*�3�v��hp�g̨r�j}[�����(��� �Z�L:%HeQa#Ef�#��\+���4�i�dW�(��do_ 3Xd��1R+�����R��^��4Ҡ$)(
C��G#�<~&���k�L)RF�{2[M��d��B��`jE�G�pjBB�i��tL�#�B��V��.Z�	-@����`d��Rk��ܨdHb�Io9̙�����
�$�����I8ˊ����?i,�[�r�������h�w��	B�0�<v�j�k= ���T;L�=��AXsm242�̼\�1�u��Ku��G�A�rU,��¡$&\\�[OGq��r������QX�J� �֦�0asJiZ�NX�L��ޫ���0��ىe0+*�-�T�j�$*ǜ��s"������
cY(��ea3qQi�i4XB���gq��oC���_a��0]�R|u�md���a�`p��/��.�p�!�;J