BZh91AY&SY��Nb �_�@yc���g߰����`�����h��4  �E1����F� �hh��j`R��h  �   T��UQaF�тbbd0� JdA2I!��h=M@`�2 �sbh0�2d��`�i���!�*I41��jxS�OQ���z����zl�	>d�T�E�I�;�Լe"SA�KOk�P��u��UU^�q$�QJ'���&4iO���/tK�n    �B � H ""� L�̏��p�>���'m:�P��(�P��`(	�	8�ܛ���Pn��]A*R�N���4�&-mܣzwT��B�%n�H�ǫI6;��]�TY�!$%�!Ho#RY�c���7.�_f˼���*t`H�yg�j�0%rb"��]z�+�kv�i�{���{���A$�I$�I%���D&�$�$�$�fbR�������������444�(�-:�n�!f����I��U�Z%{u��*����5��|(VI$����Ɍea�;b`zD�X�T�ҥ��]?��t�ޱ��J��m���	8�ȹA�4aAu�R��T��K��,��m��{�qQ4����:������nVw<��r�m��PNc��U��T�BY@n�vԆVSo�Y��B!aʴ�,���0v�w��ɩea��ڬbٴ #b�֟+6�:�[m��q2n�!�g-���PSDEq��"�$L^�CF�]C񐜡�=�>ϊ�����)��1���.V�[���A1W3TJL��ЋMqw�r۵�l��m��U�^��5�£��㙒�-����X�F�"�1�i��@�kڲ�J����o/-Nol;�7�Q£X�2���$��D#�C�d`/%UUUJ+Dh�a�AVM����@����F6��l�0B]��EUD�/,:�V��k�J>]ѩO�Ԉ��IV˷��[� b" �U&j�$��V�L��*����,8$����qy[�U�*Uz*���TH�Z}yOA�h�ȳ����%��ZZV�L3`�EJ3�X��>ʖ)(���*(�zR���b�(��*QA���sq'A &�q3!"h�J�2�A0FQ7dH�!E2B(�ؽ�Q	@D	 �%��=�C?s1�� �'�
�%8�6��U��Œ�DbB:��Pe�ZC��6�R�|�fr�%-� a��t��=EH˥� ��3��e��pĄW����sO	H����a��<T������!�T�KH�y�'�dG�����dD�d��3�9.C����xP��l���!��Vg�UKKO|�[���U���^|�2���ӦaE�?���I���x�J �*$�o�b��b�˭3�����b�ǌԗ5�$��
�*P�R�����ɔ��v��f�Q����b[��r-�����r���M�5��>yߗ�g��8qe)�AI��*z7�N�i�o1�t�b�&�����kN��Tt�%e˜�Xߜ����	&��D���H¼�������Ek2t�JL���c9�Lg��~�ɉ$�M���^���&s�x�������L�g�tT�ڔ�Z�&I�LBK�����^]!Um�̈�I��SZYC�z���N��l,6���\��Nrζe9��,�'qsv᤼H��L�v�Q���ΤD�w��1����\��Z1�Fa׸�2���b��&�i�����m��&zӫ�i�ɚ��R�su�"&s��lcT��j�-���Qhpd�����4�&L�r�����-�.���㞅M9��w�f�6����+iQ���s��>yܴ���DF��'�.�p�!1���