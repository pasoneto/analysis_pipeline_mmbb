BZh91AY&SY,^� n߀@y���g߰����`�y�璘��e�
�PIi�К�(������ꁦ�ɣM�Sd&Ԧ��� h    *��������`L�4aLC 		ML�ɀi�6�� ��bdɣ	�bi�L#0I#SA11S�S�&I��=M 4��=CNH� ���P�s��a$�t�����`-�0m	P�&h����9�,�%�i,&��Z>=��s�rwz�UT�  �"H @�1DH� !%ɪs����X��ۜY�1���&m%��P��t�u#`�;ћ��b$7���;�VTD�PaM�0d���'z�˵.=����l# ���1\%E��j����Ylo7%C�j !���E �^H��	Sg��6��:�M�m��a�i&�V�i�m�nD��m�ݶ�m��6ڌ��y<�&���i�S5A��ps��ٶL>OV��D芈����^)����暠�\����	���=5�wYD�ͅE+X;�J��:ų`�cV��Rc�*s4��-�M4���i���t���b���{�,55Ek/i��*�Уl�Ωy�n��M�Z��^��0��i#ԉ���	$���ɭ��.EF�嬦�c@�ta@f�քF�p28�Z��I��َݳ���>���$�$�_Iw��uߩ��#��i�d�%�� ��imn���2!㾴5�����I$�]��e�8uG���Jъ��-0�	���|�͌��v�-�{qI$��S=Ee�cj�7�4Z�%	��Th�[%�b���0f��I$�U�]s{�7�͞s�uF�g�.���.S�p.R-F�(od�0L'��Wx�2jF�7$#�=�kU�s$�ࠥE��J0f�=�DDD��̵3%@�۴�d{Fl��Q�	�;x7l�w�p�����$�7(N�+w�P`�xv��g9����� ��i��o��lL!�s��@���򟍡P�Z1]�
9LQ����"�D��QE
�QET��QI�#p/A�D!]���QT�ZF��DS�e�!�5��;$3 ��0Q�;^����Q����������K��\���L[f|佟\���rdp��O�0�̲�1�n9��R�1��!q(��o���ya�hlR"RвzS-S¾����s��t���X{8w5�Q��i0,\�8�Vnը�0�u�\V�a�;IL��
��λ��������:�jzz/��/����Ie1 �N�Q5�.Ա�y�WOb���h.��e�
�$T�V�e��|�vO�t3�SCt�)�]nsc�z������,R"`�,f`���u����éu8d�b�y)��N9s|���K�����fߨ���4�����.��p4F�H�z"y�҆���;ر¦��ui���)5������T�ft��J��3ޝ�Y��T� 1�F��VA�;��3�֥CR����z��D�\U�ߟ��V�kDNl�`�N0��hD=�faD���iˬ���Ur�+ЛݶE���c6�L�Y),�<ҥN.�Z"t���:�V�;X���S)�UIE�C&�o>.f�oD��x�PbN��q��2B���BM�%��wcie�b���e��L�Ȼ�T�v��hw�������ĭA����Fn����v�3,�vu��!��:I�_�w$S�	����