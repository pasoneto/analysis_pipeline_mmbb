BZh91AY&SY���| �߀Py���g߰����`
�������   a�/��ӡ���S1O)�FS� �4   jz�A$      )窠        ��4$�=# �P� @ U3S@ h      I @J~i)�5O&��=OP�2h�4�U��:�DL@�$̅"-�0���r'�l`^Eȣ`|��2.Q]�"������9C��vΖͼj������(��v՚VQ�  ��  @  Q��U�8$��+�FNJ�$���E؀F���y�u�0���i�E\g�F�
�q��(wf�&Za��1{Ni;�s���g9p���˽���3��?�g����>Us�7��z#�2lPn���]��(��Ƀ[U<��MPKS�i��B1y�M��>,EU+�b���Z%َ7о&��;�7���'q3fI
B�c#Y��%<!	Sz�=�{�c�E�%p�I_ �$�[w����W��|�{�W��^^BD]�L:�C��e�xG^zWw!�k�[~��0�s�ZUh���a�T���k0��i�l,��:h�A�E�X�'�b�x�2�����L�!.�n�t�DTz�v� �0ѫ�?S�{��F#P���I��cEc{8��0lx�7$; �����Ě������nɧh�9�95���09&2�(��SH�hR^��U��,�c����6CK9z��x  ��rc��;�e!3)�����H�D�3d���nQ{f=堚ɋ0ph�˸/v��8�w0�<�a�/nM'���Xv�nY��i`漜ڣ�{-���9~�O�}�0�I> �w'��~��jb�.m��<C�w���TF�m�Xydܐh��$�<����:��A0�K��ay�+tU�wD9p�N�(�Iy�z!�S��K
aL4�d���t�&���nB�whg���,4�6���e`9V�mSE<�{�Zf�W��A��$��w���8�y�P��Q��hF�n6t��M� �EdI��A홃r�/M�{��&.�)��F֌j�|d����y&i�$��<�x������9��N��ht��<۲VV,DZ�\#c�{Q�'+��jnJC J��d�FFārI$Զ���CE���8������L�~,��'N���,�L@����2�+y)�d�":�m�7�uc�4I%��ynx���Ym��b��D��s���M�wJi�M"'[5�����)�a6���X�8���kTT� �*xn����6V�٣����C)��|����k�"zY���R�t�������< �BN� H1Te��U.'cE��>>����(�0,[B�/B�
B$B$$_)A�҂�RR��Ղ���� h4]��Z$�YZX,�3`"h&%ʒ���v�$FA�5��R�����՘����1����'@4��O���@�y5&���x0��²?0$Ů�}-��p�L�0�0�3�2&A����	�r�V���?.AXD�"�>!HB4>��[�B�׼C����C6u*���9 ����	��vF@Y�_@��z���ZI$�E��GɢQF�J ��;L��V]7�me��Ѡ���~����ʂh`� �ڷ�Lz�m�#E�}��n��Pu��B���D)� H(��F,��r2b�B�68�mGQ���!�+�w��Pa���!�~2PDQ��(1*X��Ӈ�8�>R�I� "cx��(��5d �p%2S��
�w�m:�IV��Ɨ|�0v��lp'���04��U�{� �A�,}��zd�.�@~&�b��n#�Bh��x�1$	<H�Q�9���`h�/9�0�����÷R���#� V�Q0�inQ����ެ���{���HQ�����f��vgG�y6<c&���h����n�g$����!��p���(��
�����X��(������ETUEEV*��#EUQ��*��(��V*����/7bЈ0����#�:K�]ƀ! d���hl&5d���Z>wy�O�X�d�Hsm2�Y�v���j���țSY{.�P�0�mh@���S����dd�X��^K��mD�Sg(	�" Ѳ�0@��q�Ǘ��d�M����H�� �r׉���"�(HQ�y� 