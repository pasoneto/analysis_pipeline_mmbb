BZh91AY&SYl2(� b߀@y���g߰����`	?z�g�, d���=LA�@    � HFE h     ���z�&  0    	5I�OD=FM Ѡ  hi�i��&�&	��0`��"�M4����ŚOM=A����=3���TB*��IZ����g�`B�!�p>�Uy�Gy�	v�H������N�0H g@�Ba0�3$BC�! ����CUwwBp��3߱�}���&c��[[��9ւJf�IMz��\��u�QJVbX(c���>�� ��l���k������{EG^'w�Sv�}]�\5��V�u�su�����w}�N�֦uO��/�i&"6�RÖi�;�sG����L�@uX�����YS����c�BD^5l������X(���V�Qm+,$�i�U[V��U�Uj�\t����m�B0H�o��os��=���:=��	�oJ@P�����,�dܒ[PG��V��c�H�n��2-�%t���0����C�B��h��v��)�ܠfd��:K4�[�L�K�h�N��V�>:zK�#<˂��$Ҍq��w/�T�����C#�:(�t:LF�%M�%��<"���4fA�i��yɔ6��4oU ;�QpC��Wǁ,�5�г���yz�M� [�x�Y��:�<$k�6\��uZ��qj�~�G9kU��YC�(L����C��@w 7CX'G6�fu�u-\i���U�[]j�Z
��{C��ޢK	���"z�:�YR�{C":-��i�Q"�OM:k�&����|ݥ:���G�V�KIh.�h�y�dF�F��<�2Ǭ���l�F��Vm��эQ��3	k*�/fBQZ��]����b�Fs|C�'B�[Db/�r�4�����r��(9m��iT���h���Ѩ�����6�ݶ=���%�鑪�3h�Q�'���-�rwbݍ(�y�6oc��l�J���#IHf�L�f��ͅ���߬mp1���ﬀ�鞽|�xN���^5U@I!(��g�2�;�K4��ē�RYb�\���*>P�HD ����1�TH݁,�CV�*an��*��]�M�T&h�Fbj�J����^�Aa �BJ D :�ԫ�
�ΰ���Ȳ�,ܕ�#�5=ˬ�!�
��~|�����ߖp�{��Wn����=d����� �C���Eas�=���O���>��3{XP�����ü���W���S�8s�H:�>Ziآ?U��@S1�\d;� o*s��ڈ��ʔ&6�ͣ*T��n�T�D�1{��2�R:).������b�m@�CUW��Q�P )<����i�%�\~v�p֟OC��3�"K
$0):��9&+whOa�Sc�p
h���!"A�v>~ ��y="�S�D�(��)�1@;�<����@Ӥ��$�7��a�hA�P���g�j6o��{����Q���O��j���e+��D{� !M���9H�\���`P;�ٳ� l��TDlH:���>޾Pd��@Ŕ��&c��Aÿ4T�ć�@NDb���>��$�y�����"jqzTG���=�����i�~�N! m���t���'#���d�'��
��@b�T��C�C�n����X�DH�R)���

��ŋc�"�����,�@$4HoB;� �9�,� *�pJM3-'��A�N���1��1��ㆶ�p��W\���6���f	�G��v��b�Hvۍ�� �X210���o��`r���wbq���C�Aϰ�l��˙��@I3״�ܑN$�"@