BZh91AY&SYmI� ߀Py���g߰����`	_z�=鍚P ��:t4D��$���SjLd�4��@  h$&��D���      "��0&�L#hM0�4��LL��&SI ɠzA�  F� 挘� ���F	� �
�F�B�F"=Ҍ&� 4���OS^��'��"���H4�q�Z	1!��ĉg�0!D!�8�_4�DN�D�Q%	�K(�Q���U*̘Ӣ@�	 ��@;�'a �I � wpC�!�! `IИ b������B��6:ի�#���21��c��p�e���kz��qsg&�L�#1�jZVB��!�B�Cn�����4���x�Z���l(\�v-��'>ۧ��FP���DB���{�����L;M�n���;3�o�0������c79'����L�����t��j��/����s�
���i˲�^��AV�ӳC֤�5�*�����u�k�����v��`�sˌ;(�L��#C+t#��2�T2��Y5�D'Z�;�z�8�1��`AL�o�\"R�&�i��I���r�j�E�����"�`�����;+��t��MB�yU�קfǄX�Ԫ�1��ڄ;!����wt�nǣT��(�n�#�>
�]l��Ky��8ג�w��j��s��g��ʜ#�ul�P7yNKkZxL�.�oL�#��K~��뺷}E��2VM?;I��-�ڂK!v4�U$�Ӣ�E��j�	M��{���#�Hn��WZ����C����՜�%��9�`�l�b��N�[�+L��Dh2&s]l�F�8tﬢue�;V�Nhv����[�se�F�cU�+,�2d�m��pi_86o�nlU���<��;��$&�-ф�7̴�ff~L�%�.t4>�����Ls��w�6$d�����EsWʤsȎ�Sэ��\�q27��f��ri���x`(4��:ã�Α1����s7Wbt����1<TȢ��22t�1�j�vv����z��U�Ҁ�ܪX�Zn��UcM��7tx6l6#�Y�pzl;��Ob("#�UQQ"Yi���U�C�e����+<ح-+L&ѕ���jФ��%�P�L
��i��.�$�w`\���`L�Q,M�0`�T�jΞE�@�EX�j������j�?�\�-K~�n��Պ����a9Q=z�iO
֘�6%���ҹ8�M%�@���2���C�aX�,A9�g�/�FIu��D-,i���t�U,=#F�̧�׸<x�9S���n������u�h��{.�CRld�9caŽw]�kJ�*KK�9��U--;�z]7	�M�Y��E���ג�����8���w��9(A���F�"�ND��2Qe�L��vn�2Cd��R\נ��B1�1	��v����d�v�u�f�A!����!Lёl��F�Cw/&�|���"&qh�0��vN/�i�Le�)0���l�������d�.�	К~3����0i����������_��MG
���"v��o��d��aG5��Z���%����^s��p�ؘ�K�M}x��ռ��K�L��o)��`&�M��4����1�L��ĸI�ĕg�����V�DO9��6'3Y�B������}�f����ï�'�U���&e9��d�}���۬��$!*o!���L�,Qb���" �����`#`(�UU`�A�����bfHfHT�v˙ǖ]sVh�U��ihel$��&�i�s���vAp*�}���Q��h<f�ך�!
��;ǁz�2�i�e��D�Qh]౼��x�f��qU7.kfȘD�I���SN�~Lg>m֌��+�ңt�/�7d�� �Q��w$S�	Ԟ�