BZh91AY&SY��>� �߀@y���g߰����`���Ov��5�l�E4e=F�L�4�B=!�CCMG�6�M)Jz��d��a�  *��������`L�4aLC 	L�6��@d   � 昙2h�`��` ���$����O"6��&���2z��(A|J�ADK"��5����	��0�>�ȣ�|��y%��WCȈy�TC(�uup�¸b�-kZֵ"I �D I @"H� @E3w�ʓ�L)>b���YS����[�-;�eT�g�� n6d��9����_߸�S �����A���C�seT9�wW��o��<�S5a�gZʉ�r�У�hs6�"�T! +x������'��nf��YO>m]u�I\��N�H$�$RA)��I�$���T�Q
�P�$�2��$�DBYa��1�	��~���\4/��q�C�;���I$�/<\v|�SS5*��k6E�صp�s$��"$��݌���33��7��1�Q]��cu05��X,�cG��p���Y�vF�-wZA���s2�ɬS��0��Pl�d�̤��ؚ���~ ��[V�m�H��3�Y�m�۴�:�YE7����&���x�����@N��i��,Y����kb��5JJD
wD%��ޚ򙬴�m�Xf�6Tn$IZ�D�V5�;W%Pˈ�^��u�7"�Ҏ�]���@   .��&�m��v�1��F�����1�ZW}=I΋�@t@  z�m틷gv(��mYWNO1����CȚ�������    ,r�qņ�
�U�"�1VP�ܷz�y���J1m�	  ���n��Ԯ���5wh\���iJvq���̧�X[��uր��-���[��8�	�oɃ3B�X1!޲.t[Ļ���%��k��\m�����T�kI�s��r��~Fo���w㴄$�I$�4Q�����3qh�j�����z(�ȱl�a���� Ff ���R�$�!�`D�J���5�ˋX&D8�� i���Z�	Z���)#�{�;
PdTd	��
�O�S����K��9ts���4WwfoƩ���ᖼ�/o�"���	��|�H9�{��{��%°��
��螝��]f���8�BB��@���\�_�ӰN�����;ݛ�d: 4�ۺ�R(��fDd �58�VsxIf:�B��s3�V��"`�c\�7�Z���p��o�Ͽ~���y �0V6��LuV#W7�3�:>�-i��4��@�1�0W1�xd�<�j~�5�2:���m5��\���gV\�E�XxC�/k��n�0Cva����.ל�-!��r}p�l(p"W�p�A�E�`h�
���B�.wD܊<O0�6Gy�,vZ:����l,A�Y�{0`��pk��P]E`z�9}|�[!G�g2�PBi*Oy.�]�CK���#Zg*�d���\	GW��Ӵ+q̄���[����n�hu�1&�Y���Y�CdV��9��v�J=����k�����@Lc�sztQ���(�\9�����6�k�t��!�^�*|\�Z4�v�Q�-�5P�&ZW +Z��-jHV����w1!B�P��h|Y�����كA�)Qq/�MQ��oAٱVg��������
�wD��a���w$S�		�s�