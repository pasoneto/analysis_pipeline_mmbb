BZh91AY&SY��J e_�Pyc���g߰����`	y��oq�� t<` �IBOP��F�� b�h���@"D�       ���=&��hd�    
�h�   i� � 9�#� �&���0F&
�@�i�F	�4�ɨz��i�G��4�7b|{�!a��5'�;����Z�i����h~����?&~�~J��&�<0�����ŏ[%���  0�  0� `"   
�B4�d��
��U4`j'-7����챲�@v(�F!��Ta6�3��:��K`i��N��6��Mӆ����B���V���t���b>���sH�8E)3����6�V��h�d�s�U2�u�T�Ջ`�U'��~��t9�2���,�iϐ�q��9��� �A~O۫�xxw���33wYwsw#0�fd���L�E^b�ř�3S33Y�s33&f*�q)��xh4A�?g�}=K����2V�����tN���NqE�ӓ���� U�[8�hz������S�Ş�#j�m�Ċ51t)Xg	��p#��`5=�F�d����`"�S�ٳ1���ծ4+�r��� �+�� �-��� �����kD����e�
{f��|=Ɔ��Dv�ݡ�#�p�A �v�G�Y{$�dwEq�F
x��U�T��5���r+8� �)&ap����s��4�L��;hV�jEvA �GTc���T�;����@����9��UF�06��3°�ޓM�Pj�CCR)�9o�nN��H$0(ꠂ"﫣��*o(QAa|&4�V�L٨��*��Ps	�Ԇ�Z������A ����)��c��-/	3\5UXV�Tq�ͺ��R2�S��j��A�O8�I-p	�u�	�p��K��&�n�o[���A��$\�H���ªh��(@	�H}Z�����vS�ag#,��b�-�}˜�yxj�`Ói��y�f�$�vX�j�o�3K�nk���F�Kb��9���v}�x����:�H9�������@�]�`�3vS�C�%93�E����[�:�G����h� �[�U�;�����6���q��ڶ�W.V�L4i���]"��.P�<V ��I"fÀ�	��09��a���C+b9��C.q�r� v�Vp9#m�F���I�;G!�B��)��E݌n�����|���41�Y�e�-�j���O|�8MP�����iP���9l��M�_JyF�( q0Ø(9L�1�B�q����a���Q�a-u���6O	P���RǴi��S���z�1��1�r>E�xO�N؏�����~�D�d˭��ɹ�Y�cc�����jR�R\���Cᮥ˟�j���pa*ҼZi�f�S���W��L��W�S���Sy(�YPJ0��T��3Ql�5|-���d���z���ۢ.T�T�R�J*�4����5I��_��H�<�Ⱥ9�L!MC2��E�{�5ֆ9o�*0�%ǚ�	;������{S�S9Og-rQ>4�,Y(�dU+��(��)�b�����5�MRVq���+�<���q�$���o�*F����
7�&�l3p0�7����M�&S����ΙH��sx�3�{x�،�M�b�.]W�V$�פCa��O5�MR��=锒%�IV��u��B��NP����6%�}{���u���X���Չ˕J����i-���p�`H�0k��QGc����!@PPR����IIUUUUEEUUUE	A�9�4�^s3\v�M��3C���2��ek9L/�γ����j�4؝�����s&'c����IМ���]�]N��;���۰;�T�5�l炩����.'�1I���tP��i;�'4Ѿ�&�.K>|R���i�kx����)$[y�.�p� uҔ