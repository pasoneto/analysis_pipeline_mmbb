BZh91AY&SY�o�4 _߀@y���g߰����`	_z��J��( ��P �JjI��S�<iM4��4ѠѠh=@J $��LQ�	� C G�UM�h ��   &�*Ch�#L���14�4�12dф�14�&�I&�ɒd=��S�yA��yO�����
�uP2�s(p����g�`B�!�`}���&��Dt	���DCǻ��w�cqv�[Z��ջ��.����  �   ��	0HL���+�2���g���~
Ο���#
��n��كa���6�$0c�A�\ f"D��.�&i�[�p�==Ăߡ�������,�U�J�'��zYU*+M֕�i��ʝ��Ɗ���U�UUUi�j�G�B�B��B����<�z�me@*�3� ��;zb?��r�a�:eUUX�USWJ�WJ�j�ͨ���UU4�g*���U�0���P-�u�5��$$H0�?�����Y>q۪p�|�<G��D��T�y1
H���Kf`�A�򰇣�9��H6�L	Av���,2$�*�?�}�;��,D�nFp}�-7cF!�@�!+$u"�\`{k�ں���w���]Dh�lA�&2�.p&c+���Ƃ�)�&��ht�t���|!7b:��M0�v��yW1�J��L�z��JR�7���^��$7��:��آ���b��K㡰��A�X�u�&������6�x
!}.v�G]�M-�b/��X��!���='m�0\qQ#�l�V�s�"uд�����Ĵ�;>����#1�A߀����*�A�X�����,HC"9X̃���)�ZL��̀֫�W|��A��{��m����\V�k��u�(1`tIw� pФ6��i��CM�֌�]��"TLeA�����ܭ5�1��E\�H��=e��9b;9�|*���'VM�a5�ۈd���(2�����5���	\�[韍�s�4J���l���$ֆFT�)ڶ�ɛ5�ȑH.��3��5g	@�"��I�|#�;%-!XĩBF�'BJ&;��No��y�"1{ꪀ�IEM��@h�v�����y`SL��f�+b��
SeZQ
�P2KYdE�A,��]2�%�@���vP;Qn�����:���b�H� HH�٩�L���3D��~�yjV�����4���hHF�<L��6)�()~�4��+V��TF1M$�QZsd"*$1�+�',I!b�s-Z�f�]mW���)@| �hy��l���@r�	�5X���ׅ	
�VG"j;����
��ҿ����#M��i����� Y�3�e����=�p�<[@���y�7�^��� w�_PAF��J��&�b@��NJ;��d��S���n�)����`@�FX��'rf�;½��Mξ��*�`Yf&!X�O�V���|�fa�<�"��!I�R�{�zc��^�˰��(�r��������=��.���z�O��_���EF�d�����pC�iWS�|����<%�u]t&���,�7��K�z�����8#r��� 2l}�OX`S,��!�S�k q��E6�#�@�C6T\G�7PZ e��v�� IX��Q����w��c!����@�ƤO�ot^�:p��<���(Z>/�`����E:&�⟩�1błŉD���1DbE"@�����DD�#�����ѹp٘�� �AHcVXP�ڹ��<�_��3����s�k�� ����QG'�7���
�y8�7��`R u�����n��K��f ��qo��C|:l�w�Vg:LMy�N%���?�3��{X=��]��BC1���