BZh91AY&SY�� 	�_�Py���g߰����`y�=:yD�{e(�@}񾤔*[pZ(ID�MO�"4�hdѠ   %O@�����d �   ����f��        4�UDɡ� �      E"hD��SI����z�F� �MD�!S�4ɲ�MFF� h ���}GĂ1��D�>�l{��ؒNV���kxdl�j'h5$�L�M|%�o�6����X�P B�����mݲY�m�t�Ns�撀��� ) �*� &@))Ϳ�8d��O���Q�s�"_�$�ȹ���.�h0.A��<��sOJ��v�"]��檖��K��j{�*�����O��M9�
"]F*�}��A��|>2`^�|�+����}�����s.��}�-Z�_�krjd:�,�!�d���j������M9�
%Σjln{J�.$������#kO��sЭ1E-�BB�I�L`�C�%����Bv9��f�����NffF]UTϩ�n�����n�����S����ܼY���3uU��337/1[m�⮔�)l8e3*�$F��\���qO¹����|��G���|^��dA��jҊ�ȃ%=ځp��$�gc&L�9�`�Y1O	M�>����sf�<:4ݻ��8V��;�l��o�q��mߜ�l�<���*$�d�ffL�0�ɃM��L7UV�<��U^O&&���5,{���,t�˿kp�U��k34�KU\9V'-1�D������OQ���wF����cov������&�fffM�&L�*|$�@��8��r�ݦ6��8rƕ+�*r�
�]k��ٱҹi���t��uiN�Tn���f;���ೲ��»,l���<�<w�����UUUZ9�/.�����0��慄���t���a�1&�0!�$��A�,�	, c���4�}t��Ɋ�,�l���ݫ-��5J�����j��l\�b�gv's���n����Ӗ6�M�O �d�Q���$�x0�Ό�C�:A%�Xy�md����������<�4��S[[�N��\h�^�J�v �`��(�b�a�Qe�d�PBz���A	��#ֳ3335Ba�(��^%n��c��^t����fvt�]0��9�:A�K4s�(��'�/.f�L�2�(fffff�It�ic�縣M0�xш GK����ệN����r�tݺ����q;�(���3$����A�|#��a�ڈ����ĥ�'G$Fb]$���atЇT��M*z��;sIr��
;IP�q��EY0�A%��%l�L�财�BG���Y�0sDA$���p>����%U���im��%ş�y�Gσ��1�Y��|�|�2d�q��G;a�\��0����׭K,Qe3&&`�K&VR��������2�L1���Q��bkZ4�Sj�ڦ&��I��Y���%Wif�Ȕ����r�$��(�K���X«[�ylY[��-�M��9�_Ј�ţ�"�>�Đ��5L�`԰G/���Ɠ�,XE���Ee��aefŦrc���I�����Dd�����*ٔ�'�LIK0|��[?#Ǹ'ø0�%:B���*?�<�ص�{�"wO7$�����7|��q����c!.jm�2d���0�%I�!�E�b�ek$%D\L�&��$��x��׶������)��`���'��S�u���OW�Ӆ��>�\���d�X��```b%�e���6-n`��)��<f�Q�'2� T���>�"D����)����F�3t��DLMN�e}Yԅ�J0o-�"a��9x��o
>D*B�G����*��At@�aA.�8VF���	� � �T|GaK��n�#T�o'Sҙ���JG���f�y�4sO>T*VɒL���ˠ&!#�P8�5VL�T͐���BOߥ�*�쮦e���a��a���OW���=�H�`��&�(�I�9���ϰ`��E4��@NP@�1�j��F?T����l��ww�>4R��}��|f�        @                 !�$Ԗ��0jUJT����/ʜ#�|sdxt���,�{e�LL(�udJ�ZB�m(��X*Ou
F�!�|�����$Ng�p���U˙��N<�hy����h��4>gS�|\J٘�;�C$��������n�?\j��%�m��3�
./����1��ܖJQH��/�.�p�!�rJ