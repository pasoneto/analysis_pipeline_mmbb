BZh91AY&SY{�m� ^߀@y���g߰����`���K@�U����I!4h�ѧ�j�?Rhbd��h��L E6&O�Q @    �ߪ�a4hhт0��ɐ2L�I"���   � 9�&L�0�&&��!�0# �!	4چ���!�hz�����JU(� `;�OqeQ�Ǹa�.|�-�F9G���w�D]�W"!��GIٻ��Y�~�Z�ikZְ	�"@H�L �$� $ �'Ο �������"(&"�'�_��M2�*@.��vz5�R^�X�K:�)/f���E[+Q��ڐ�Vh������L�󶔾:.�����sT�D<v����J�����GUH4�h���]��v3�h�)W"R�O{�$ * �(�VJ�
 ��@ �   ��-�1b��	r\�R� �g��gsٞ��]σ�������Y �e�Jv�9�OD#��r��$��KKd����S̋� ��;0��� {e�5$�A)v���6\vL�vP�g%3�QL�
>8Gg�an���l��2`ۋL���[�Gi���^(�{o\%I$�JGBs���#��yP2V���a���WH
"�����H�0�ޞ��B�S��1��1�`�I$�G���w�f+�����)�x��rŜ��;A,��' �a-��I$�/euӾm�.g+*eS�MDf���/�興��3���I$��;4v�*��a��+��T.Ƨ%ҡ�R�!�˚�bI$�V���=�((*�+_�J���f�n���f^򫑁�"�&�by�y٫1-Z�)4�h��M�"��k��W��fS��O�I2%��.\�GX.ݱ���'n�f9�����������I �s�$��S��sq�`�{��%�x[um�C�$D߸Q�$a!	=rI�|0y���0Z��~��KdX�`` E�H�{�9PS0#*	A!�( @��� ���KT[Z�`���
�( T��A4���B����Q�x�ddI���\7���GĲ����q����-.��}�[f��c�Zp]?\K{�uɃ���v(�.0�] r���B���Dz\w������ϝ�vD�({G=����]���"a�j���1�G])����1�i�52
z��xK�����I"QN�+o�HA�f����.����4�t<�Ѡ���Ƈ݋?H]|�9ثV��;����=��O��e��ch]���
�F J�3�������NVGa���1�[�N��~ݝwe��A���eR��y��W�SaP�+`�F8�����2TQ\� �3/6"�N���B�Ml��J����X(��#�zF���X�u�hN#��qg����������V��a��۽�w��(#6�?R��^m��Ɛ���4*�dX`Ti.����ټgP�B �fhV�/�ea�̡4�h�뜼�ȭ[xtg`�%����5��pQ��:�ǜ����%�Q;9�Qwg $sSëK�Y#8R��G������,���#2�iݒ��*�%��h�o5R48#���dff<d�&��>�!�M^�b�Po�@�a���b���L���<����n���)���mp