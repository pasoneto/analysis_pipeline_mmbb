BZh91AY&SYS��$ �_�@y���g߰����`?{��:�T�r5� :dD�CT���?T�@  �=M 5OL�J�MM  �   ������  �     �!1�Sh�@h   �MS�@ Ѡ     $@A56Be7���?D�=L#A�4yM��-�� ���1>-���a���[/�F+~��'΢K�%4�S<*�ϋD��
F�RL�ک=�^��M�G�64�]��fX@
�  � ) �J� K�\U���J<�Q3��é���Fi�3���Fj%�F�V��.K�NM���][�|\�1�XM�Ua�Ea�!UP{A�����$Wul�+��a+�x��p����taeֻ=�q�cz�\H1���c�.�I>���^�;������@P�("& D�	 �D@P� � " �+�����e�l�2n�&8�ip�\��F�����ΡxA]�x����I%�6���l�s:�SO"�ƝT5��N��(H���G@X��=�ͧI$�J��b�H�%؃�&���`�K$��r��ہ�r�bXY��:��MDǀ2�f֍t�?I�uM�]�$�J��p�{Hc l�*�)���E��	.b��PXI���5�"]A��裼U��%��B�2��~@��X�I$�,��4z쫳}	z&��'����{��Y���x�n�t1�-�Xܤ�I$�GT��a��[�茡3��/CU�E�B�d ��{�;�Z�Li$�I@���5pEu�?[��u�bn-��5#Pq�t��51�zS��0ՍĒI$�jw�r�\����|9�jukM5�x͙Bl�T�4�;;�>!T\Y9Z�U�g��䙵f�U�RV31���P5�$�x�[ѭ�k\��ǒl&��)�h�b�g+{�YfL��lb�>�Rb�"f��v;�L�px��7�]���%�[���KH ���Hb�5�}ؽs�c?)f+��p�ʾK���b�(�E=��J*QE(�YR-(��b���*(�����Zˁ� :!�4;��Y9� �NB ���#Ja�����ab�S*���K	� �B 2����yb߂0����������~����51���c�*m:�F]B.e�y@������_Eٷ�	���4����շ�}0�lsQ"|e�d��{��a�m܎�S�R��N���`~\��y"}#�{�O.�'p�����&����!���)�8(�l��gsO��)OfU��r^��ϳ�y��h 8�Bx��X(�2�`�EH9$QFŏ�ɡ��"E��B�[���a�nf���=x�۵��K6˥3LV�pxK|<{s���(�.�,ej�w;ެ�9���:ة�4�,$r����zv���y����_��;D�v����>�&*��ϥ��#��cBIđ<_jPƻ]�oS�1��L�WRloa;��&NLY߆��$���aw�ό�~���E�Vժ����^[6�T�Jy*[U4Z����`*��g��*���H�j�;l�R}^�����w����qï����ج��K�i+T��,�?'��tmM$�MG5*T��u���D�'�lZY_�u���5������d�p*L�!KM��/3ѿ�zis=���L�3a��zXe��dH��:��k*Ζ]
t�K�*�fk��V�Z���N�[X����F�t�IM6D磜��Փ��[ԭ�]v�.�j��T����P��d�5ɿ�ܑN$��� 