BZh91AY&SY�䭮 �߀@y���g߰����`
�z�y����� �s  0!	H��j��jdi�`C&�!��5<���"��@   4 T�O�U d�d1�F�2h�@h�MH&�)���5��@ �� sFLL LFi�#ɀFI !��L�G���M=G�=@����jk�u�
���H'�s?��I�A/:�:b.b($#2��O���	&�A��$�TYHƦ��vwu��w_��	L M  &�L$ &�D��b@	-kZ���M�,;�V������ޱ�_`�y���ʁ3>��}<�ɨ@A��u��������혡<m5�y&f�a(��dS�!|ڡT��>�-D�-�Nb8�s&��4����ԙ���]ɵD�Q!�7(�t"\�U����M�q%��#�n!�<�k�=o!��Su��=�4�I�ͮ�~�{�������-���wuw�[���-���o-�;����n[�wv��9���cƷv6�m���������;C���`?��z�������d|ta�2��\��Duki3`�w80m�s�G���2s�D�0�����9�B^��&�Dѣj��m\a�~P/�89�\x�܆)�%�]��@��El�G�}* �ׅE�����\䠻2&���1`� �8�ΐ�5n����3�� x̐M%��a���!q��D�\��b؃�:;�5����3L�x'XI~^y:�n0U�*�$KKχ~G����I%�{lpP���%6�Z\g4m\ڬL%�N�,��2�	��-��lذ���U)�6�,�l;��Wb3�L	��T���EW0���D��!WLsr�{��3ɏ�S䊣^}��)$�H\@��� dh��n1�W
���@�ǧ���b�,��$^����t��[޼b��g���7�	ݎ�	uOh��-$�Iv�'cw$i'�Ҭ�Ym�)���!��U"f1�c����������MqFM���1=��x��VQ�{�cI$�_RG���F��c�T�.�-�EėG/`WV�	�C��=�$=�z��7T����ڙ�UU���I�t��asȺ�܅-��P"��$�Y܃$�ؚ��&N�ne�����몪�H$�"��/7�y����p��Y���xe,��sA���}���!؈��Ɋ�wEwf�eۑݞ�=M�j��t�T>�'�'X<���7�bC�t<P���0�����^(]��e#Cp9"�NȠ���t��xGz-�T\���22�sA��`���o��e�b�ttX�[(�|���ޡ�8�^y~ ���|o��wƪȒBQS��y�3�Z�>~k=x,���u��1F�m@P2 ��h2 ��2��T�	DDF0���V
���-k�L
���bȵdذM2"n&�
#0�A�d�"��<�W'��ߦ���$���T��6O��Đ4zP!���	I��͞�H��m�]U�סs���!S(�E��VzTɹ�H��'�����=�>�}&�z���,�'���*a�l�Iيr)xX}&.�ߪ�P|���'�qe�D֛٥��������3�),���h~�t�ϣMNX���]��կ<\#ұ��/g:�,g�|�����ڦI;�@�IR��J��}�T��~?z�2P��?O�1�;�Z�B�
�J-ɞ�'a�d�-��a��S�"r��v�t���l���[X��<{ZL2�H�t2Z�;��~_?����S�b�,	ƞ\'I��ug�a�\cW�w���8�%ڝEe)�[�s̕��$�8�$�I�y�C�v<%ޥ�o�4V���yCqy�}رs��ߛt`BJ��M�/���]|إ�)�j�-�2��H�tT�QmJh��2=�Z{�b��������ܝ$��\w���e'�{�Y��ɴ�ݵ��݉��[�'[IO��,�O	y��5.I�@�!�t>3��UTUQTQTX�(�(�(��"���*�,DQb�,QE�(�UE�(�E(��E�L��G B B&�|2ô�s�0,ؓ�Od�Zx�WO
�Ö-���=g�{L��a�0��l�2$L���n5L��f[�Ѽ�d�S��vd͜b�`�����ƥI�LI����sRS^�O	�n�M�#g'J��ɍ*8L2��z�lH��;���)�'%mp