BZh91AY&SY���g �_�@y���g߰����`?y�  �IR�(D	���hЉ���h4h�@� �M�=O�U�&�M2b4�!�Ѧ@Њ����� �     2"�       i��&�&	��0`��"I4 %=���yO)�<MLOP4G�ɒ��T(�d@.F��y.�%
���^�2�b|"-�F9�@e���#Q�SȆ�/tD3��Ǥ64�]���.�   R@
*@ R@ RI�$J3zۖU�*��yĢf,���V�LFC׫�.Z=w��"�����b��7q;Y�W�
�(Y%䇣9��[�JR0�ʳ�4f~|#Z�	��W�@��&�0�t[	t%c@�`! $�)��#rJi�}�h٩S�[���� �#�	 @ ffaH&   B��   �iAc�QUrs��������./�=�v*Ǧ�V���#d�$BQk���fff~[��cACf��Br�̷"���JA�榨x�Tc�#�����P�@{��i$�Ix8i>���t�akb��~9,(�x��!���"��%��}���XuH��t�T-<�����30i�]����JI$UJ�����q0�L �E��&�����d�1��cDc��������o��/��:��`�8�����@w8�I$�'�o&�:us�f����m���|�{��g��5��Q�`%mĒI$����EuYY��׵�~=-|�[0/�<�ܷ2��tf�� �4�I$�zY�/v�f�A�\]v�urc5���jǧ�'3�1�Ƙt�I$�`��<�qF��H�\�V�ǹPy��(���wGI"�LY���O�ͼj��f0r�nfm=C��ΛI�ӝ<�.�:��E$NeM��r8�f��1��L��4 �N��2QpbrØp�PI$�P�m�e拑�{~�>W:���YG��q��^���A,A �~I!��E��o}]M-V|�k�
(�ıl���PP@��P@��fPJH*PA�H D�L-`���KkX,ʃMi#A
��3��Zh!���z�\
YRA$~P�D��׫<�<����vi�|?k�������ۂ��y�ݎK��5��՗ps����h����{ ���3;��ı����<�?��f���n�����!!v�@��.v���8�=�,���� ?m���~)~C-!��)��C�����u%HD���9>���3:�$�P����o�.��8UM�A�d8h�{����~P�P�A��r��x�{(��0Ԟ��0�ъ�L# � gȥ��D`P��ZN�1-b)�9e1AH~'���N��Rp���s���{��)r���u�yOF���n��p�֊��ij�5�!@��04����ט�Ȥ��� ��Q�;y�t:m+�d��n,A�l0~sՉ�������V��,]�P9�&(+�Ma��<PO����Q�C2�&!�@Z\ �s�xwnJ�r"�aa�6:Z ��fA��t��� ;;�16mc�P�5E��8�=G�¸�Ta�r�}/���?0�Y3hn��QU��
�&3)�H�D�Q��Me��ͫ-{}�B�K�v%�������Ʀ��G��y�U(�1�ChH�nGs�a�gqR�C�f2�bH�����,XL]z���F��1PC�{~3�2ԣ6*v^p�����rE8P����g