BZh91AY&SY�R �_�Py���g߰����`�z�<���mP ̜`
�@I&�M5��M��4z�P4 @h�*��� ba  CC`�檧�i�F4�2 hh� ��Q�A�@hz� @ 9�&& &#4���d�#Q	�@�&���=&�� A�7���Z������PL� ���G�Qq$ߏ�6?bI�I�e!�>�VCȪ�� �@�
��	$)xs�~�j�EI�� � P���#D
!� i�6m�@)v���	Ҕ�肷E�t���l��u�Kհ�G`dw���7hѫQ�d��Fɉ����s���#].T.m�Ӌ�;�����o�ҹ������32�br��.��p�	Gep�aC(�]�C�Cw�R2�|YA�)�ܔ��g�"����1V߶o�Z���Re�"���ֵSY˚�UoeQ\aV���Pa��n�>L&/�ʲ5D�ge=��Rz�z�s��'��Ȯ�r�]̧��i\����QLw�ܦ��73/ �CPU2��:7���$���
k��C�X�M)9h�I4Z��Q�J�)��D��1dXjT� Bj����I�A���%i  �eދ��S=�m��L"n �͜o��cF��R��g@���"�����p�e �+�-�٪��i�6�"і�13�m#X�StW�*�r; J�d^&UU�h-��b��2S�$X�[�.�D��	�ԣ�w(g��h��r�m���/�Rue暴�lg�N# �Ή 0��'��r�
�A������\�|˖���dȁ2r\ ��풺���d��gfVR/*bl��t��L�.��h�m�1bP�f��*.���[+3��A�m?PC�cE^��q�yW�LY8c��&AeI���#�������#�w�ԃ%$�W�gf���q�e[ |���IȰ�F��8\�RR�F0Ɇl������2J�XAς*fv�5�j���M`o�on'|�""/�Ȅ���w7Pl��0Z�>����$�)u �BZ1ZB���&�R�4�d
R�\�3HP��`^�K
e$&Ԃ&�X�D��k�x
!  �o�ފ�<5��ն��m�D٩,׷��$4v?O�$�	Ԁ�5�U��sy@�x�_yY��"�������i�p�"�R��2p��*�!�NS`Y7i��!X�$�q�2e#���x�����H(�������;?8��#ȷ1P�v2Y}�<�"�|�څ�INEp�� �O#�v%Z!�=/�>2�R8�uP�c�\Mh�!�
��!%��X|CjdC%�L{d�ƥ�Cd���Ν%!V�����C�0�8�=�C_X�j�;6j0H�QP����a�[qI�C��|���j_���`�=xK��J��F�Z0br��m]�L��2��؎�+qN��� +�D~C���<	=!�d��'V�0�o
=u�B�
q�ā��Tn�<z�)'�,8*ܠCd��MT���	�[;Bh��x�����4p�����X��,"?(PN���jй#c��q�t���0aɖ�@#��D�QRcr���j�7(I#&�Ha;N���ސT�E"�A0H0@E
(��(�"ÖK��P��A��&��d�")$�����f�)<��x�v}ۇK�m�2ع\���+���B#s����Y"fN�-�� ���ٗ��*?��#�r,�2R�|#o�pN00�M6W�c�R�4�;	nE����/��w�0�5����"�(HF�� 