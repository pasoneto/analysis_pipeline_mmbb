BZh91AY&SY)e&� ߀@y���g߰����`��@  {��  ր�=bde=L� �@F���dH��     h S���TCM�ha4`# ѐa���@       sLL�4a0LM0	�C`F �"2$�S�&�Sё��oS&����'HB�#��z?':�&)�k��E�/��,����|�p��=$I�T�%B<�]Pʦ����߹�c��@ "H"H D� �    9���2�64��T��0v�,ŝ�_מ݌��� I�a
#0��N*T-kle�|53n��2�:��h��$$d��I^���L�%$�!M0��^W�x��8����`�B��-�E�@����n�@ff`2�7�0��D2��y9��n�!^������s337sF���DF��ř�{���wfb.u�̌�ݝ�݈��������<�`��U���v�[��\3*Q(a�ؔ�br��c�E��h� (&7�oCy>w2��k�Ƕ�b����R���>0;�ݘa�H�$�,;��&�]'.��9(J
��w�saӮ囚�s��/wSaa����"�V�������79ߝT�Ʈf���H�A ��r ��d�Txg5ή%��q�}���62�:�nD�D�;�h"`�N�eN��6v�\;HR9:�0e[��ּ�p�	��\v�ˣ5<"��Uk���E����.����My�x�������*��@\����s}]LF��A0��P�s,7)޺E��
'��T�lZ*a�ݍzǑ|��$	�1�YWIt��RP��Ux��(
��d�O)FَU�;6l��MD9\8��u�A �M�4S�g��;*��A�d#ʱt�<D���V��/D��s>:��#TBT�H$��\��o�4�ڽ$O]����X��#j-`}%h���/k�!�1�y&$Ƹf��9�Ƿ����`��9�b1e���v��b��ҫ ��0�X��k��5�ˋţA9yf�����>��]��w~�ȏ\gD���QBZ ����ޯ)��Y��w��Y��*�_4c(�EE(��X���R�E)FR�X�e�#Ɗ���ԋ^�i/{���"в��uKIB�Ҙeh���������\�ARB�M��5�_���b�$����/�rg�HH�;j�ﬀ��$�Yv
Ҏ�+��'E�i��!LC�Jf�S�y�=�n�2nz�D왿�s���k����;"�ZOjg�x)����8�K���su|��ӏ��"'�9�;N�mNF�i߅�T��o���*K-80�9��K,�i�ъ�.���=z��s��&*�88T�����/>�0��j'D��R���;���*Y��=�����L���>^a�ۜ����AR��l���3���u񹫸e�lz�f	MI�}�	m���r��E�����sֵ^N׋�/�g�z�X�tg%FXH觟�u�>���3k�j��x5�I�S������b�p�c��8ԑ'=�rP���Y�^�&1���'�M��[ߋ)I�}�7BB��˦__���,��R�F˖R�U~��z�D6F:*x���4Z�y�Ii0gg���p%U���D�����6R}O������s�5.�����
�nIwKIO�봋?t�kL׉��R����]��UB�RJ��Q�      @  U%W*w�������q���h *�h�<hȐgAQfKGkX�%0�]��%t$�t�i�3sF9�N���H���\��f6�Zͬ����,��t�'^Lٝ�)T�bjcC��F�l�IM5��o��ыW�τƕ��::�:ԕ#M�����)�K)5X