BZh91AY&SYM�Uj �߀@y���g߰����`=�罛�� ���B���Q ��jm5OQ���=@�����QJ       e??�TL�10LF�&�2h�ѐa! ����I�='�ѵ&#1=FL�&MLL`��*I ��� �=M6��4i��A�ih$�$��"0 \�\�[$��c������g���Q&$�M{��UP�,��4����h0֏�������( � ( 	   @Et]^tS���tc��f3m̶H��0��F8���[z�˾c�fS�l˨��5���Yh��X�1B9G-��[=ӫw����)�ap�la)=�KH�8a")�1<m����c��^ڙ�#d�Җ���u���݆�}�R��Q3(%I$���������E$�	$�I;���	$�I$����.d_}#�EEo�;r��D�s)0U��q�G�U��nk���L�Ѷۚ�Y54�/�0�?1uM>iB؈�h/U"�M\����	m�u݁�0���I�,�|5�[F���8�pn�t��bۃ�P�a0�T�֋aΛ`�ۇ�����%�x~6�$,e��)k֋��fI�N3~��q�hag��f�6�;��4����0[n?Y�����y�9
|9��4GC�6uI$�� �9R� nG��Y�nA�����C��a2���ps2wZ��I$�L	���1O�1�v�p���ċy���J�����.�a$�I��;��`ʮVw
n�����3�j�TLX��ڨ�P�2I$�M���v��ǁ�DLM��cL��J&j0U=;��IbX�8�UY�b� D��W��3Ce�ݳh��;��6n�'ި]����Jp^���S�J��Ro6�M�ž�E��U���mUN���ũ���'��-�aO�2�Z�yn��oU�㻬i��lpza��lc�m�1$(C�sĻ g�B�J?�� ��.�3-0`����QETQR��Yj��40h`����C��(/e)�#,���b�%2	і�E=FZ�"�^#nrbM�$6..�M���fv��7Z��u\^i�����C�]��A���k���5���P�O�L�
eaMq�"�^q���b�lr$O��~z;��~��Kj������L�����׽�|�ɀ�f��N��q����&/��t4k73-;�l����v��RB.2����4��^!P�>�9�vw����]ڡ�SP3�x��/�,-Gy0I����9v��g��(���G��j.�@H��T�R���Ϩ�.�-�x�h�*��*�3"�:��R��_+���G*���<N�^_�����u8�b��8���9:�:g	y�b\�q��_^\5�I����>[��|wN&��BI��;�T���o��*m�hV��{&���]v��pݩ��"L	�B�ϳ����-{�`Րeݬ�/��ʖҦ�T|ZA�Ih��:��^n�U[�a"yX'cl�,�����OaX9&��3g���e�e��c6� �I�#G�MY��,�;%J�N^gI"s���]��:WYGIe��.6�����T�e���wJ�=���9�{6&��9w4籡�|��J��uL�7;se��qe��6�Y.��Y<�S2��S}�W���b�&ɶ��5C�N��v�E��\z-=�oU7�r��v�xԔ�Q3��.�p� �ڪ�