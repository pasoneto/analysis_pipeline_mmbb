BZh91AY&SYg&�� g߀@y���g߰����`����9>� �.}f�h͆I52	���d�h4���@Sh)Jz�@d��a�  *�����b����ɈɄA�%2M&� @    ����42a�4��h   $H ��L����6���H�d�R ]dP � 3�ܙ�Hf�9�|�gѡ)$!5V���M�y1!,ITh90���^����ۢ}17)JR%)d	��L�"@!0&@����	�Vuud�&|�"ET��8D��.9�������ˋ����0D۹g��j�|��C2e=�b�0�#j�&�CbȮ`���op?lɅL�0Թ��AD�2	ؿ<����a�����`]�����Q���P�:��<�k�`���N�d��$�"e�JRE$�K$IT��I'T�T�H���x<���00ط���+���@�Ő�����Yt����'h`�<a"������i�z���14eIw���7�6�#=`)顳�i��j�m��6pJmۺ�HF���z�y�&L �aL��&��DR"�e�8M�"n�[jز�`�L�~Y<��5శ�bKf��:��ɶ�m�����E-)��,Z,񜄨uRA��͂Z,+7:iV�����Y�H�vE��%"���Y���A��Yψ�]��m�����U'��35�g�.��t_�z����^W`��T.̓���2I$�LS�S�K��65��c�"���`TL\f7���V���u&�I$���e�v~��v_��� �*ֲ��o�6@��tiN�1�I$���jD��|�t�T�"]s..xsU����AB��#Ek,KU&�^yeff����ݡ;OB�P�q�g0h��]��ffh���cE�l����ڇi㌷��-��39%=333Vೕ��m�C�.(2I��Z
؟[Tm��18��9Ci��o�m�4$( �P�.Pu�Q.c��|vcܒpBI���`�B!���

( @�!ʐSh�3! �!��"C40P"u�I�2s��5F��[���M���H߽n�|߃�G�.�&��m�V�k�۴�'MU��]>U|�Ԧ&�N�&qY��� s��1h��8[���½��l�$(��BQOJ�iy�`#�q�$@�6(a�� �i�q��_TSq~Ab���2g/����-�n^����R�]vݴ5W�9J��(h5Σ4��AJ.8Ap0+��XMij&t/�x9��I[#��2	��	�H`4�n.�
���F��B�����HL�T#acʢg���%�u���#�@V��d1Mܧ�#Y`b3��iR"�[ʳ��H_QU_�L(Kі'Uv���bllC뭙��x,�aQn��Cx`���R��E��T�$1hIt��5T--Z�$�q����I��E5O"ĉ��fA�����^D4T;B�$(D�px��f�	��*HB�$"ڡ8a��f"%��[�<�i�\R_zm�@�p�jUAq��T(�d,0�/e/����IQ:�Ͱ�JV�A�rG=�%X�x���lֽ�����/�e���u˝U!
�Qc:9�6��`,5����T��(q9�`Q �?Q��/������t"�;wB��F��ky�`7F}3���"�(H3�q��