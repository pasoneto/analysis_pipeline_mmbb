BZh91AY&SYC��f q߀@y���g߰����`���zb(�'�BJBI
zjbjm=F�Q���zOQ���dѦ�P�@��Q4�h@  � ?o�U42d�FLMF�d�d�D Jz���    4�ɓF�� �0F`$����<�P�`�4h���di@Ԋ D���C�Xn�0�~����Qc��	%�����D=*!�s��{8�Ƹܵ�kZֵ�D "		 H�D H!fn�زRu��)0��E`p�b�[�e��,�o��ԝ"ܣ"I҅�j�кB���N��̺��*�4����2�q��ϸ9 Y��{�I��-z�T��[w"47�"����P=��y���g��w��oM�3t�y��m��qM�m��m�s3��n[m�m�D1�����<���� �����fxnc8i��ڮ���9���(�ꏎfߎ/b�u߲I%e�:[�ŭ��<�U��rn*�B$�aCn��:��s��,m`�U�6�KbCrҭ/I&rel�vN����.�z�r�����!��e���E�JD$K	�Y��!��<}�!*�k��E$��k�d4�dN��ʪ&l���4{m*��E� ��������E�-QG��Smq�Mu��i��c[I�b�N�C�VE�I�����h��'T:�t���5�p�I$�#eU�8wʕ��B/���s&"3ƪ/�2+�����x�I$�\�s��/��@!5}b��2����%��J�����Wb����I$��d�r'.�[ý��*�ͺ#j]�Y2UVpa{w��%���I"�w{���3�"+��,S��no�2+�7�7t"(T+>-��E"����*OY��K8��aGT���f����Y$�¹��X��F���.Vo
�>,��\�
���^`�HBOL�A��E[��a��2'ۺ��SrI��eIAN�AH A�aU�H��`D� �(�jB�Z!�S!0�!�2P�� �w��U0p(��C^��L$0�f}�:���t�<IQe;m=Zy�x�]�v��p�HN)���Z���)�L�c�E�qm���m7�'��H�V^���f���Ohm����,�C$G��>��c�0�7	�q�{���c �	�a�!�3\J���9s`�V@��ld�%�1���w��:oHؔ��Z���9�m�F�Ѡ����3�{??O cU�i�ڼk�����,n�LtO�q�0|���0�	]]a�\����g���ol0�nV�C�����gn<�Q�jXx�3�?�����\��8)�]���1SQ^��f��U&�Π�!	�&�b�;r_w�5<"��Q��0��<e�%���2kq7 �,�=w.sninm��
�6r����ol��3���aR~��{���ø�j!�U���H��_:5ft˒�cő�R�0�����"ei��=��N�:��d��V�Wq�lPu�A��a��1���Dy�Ł�z'kw$�0uk�J}4�Ւ3[��p���U�+�RXJ5��X�X��!Pr��p1���܎���# �Ȑ�sQt)Q��{��a��=��lΊH���/��3+T#�#�0��T�ܑN$�ـ