BZh91AY&SYe�M �߀@y���g߰����`�{�2��	��4 P��P���4      S�`ԑM       )�����F@��ѐ� @ %2@HI�j��=F��  h�bdɣ	�bi�L#0IMS�Ѣi���?T�z����M��6���y$N�$�@��#y�ϑ�I�ԑl�y�顎l(DJ���ͅUY�`��+�*F �KQ3T&*�3V^DG�Cr���/� IAHID ��k�
$	)&���S�N�>��.�����]�sئ����=��q�92��.�[�q$����f@W"�A8�������_%5�tjr�w��X�T�j׭��ڻnJ����n_f�����tH2�F�4�$l�8�P����L3ٳmv��x�e��6��m�m�i&��m��m������ۧ�{b�%6�<<�M��R���Ń��u?��R��F��k��8x�=�6�gW2�M�*�[�$w
J�@z�����H���*�@������
ff����o.�`wֆ����ٞ����F���m6ڮ\�ʫ�a���H��oG�ؠ��.��"ʈ��*�b.�tpaWA��) ��spF�྽t���jT�E$�,�0�7]�/��57{]��X%U5x@�2�j��UUSYrYAT���Ub�RĘ��;:�4+te���5^�$�^0�u��u>>��R�61��8�|ct�ɓN�5���J�NF��[I$�]�;���Wz�2m���u�%���5���|�putyѺ�4�E"�c��''u���HJy�7�be�-J��	c����ՒL%t2P�Wf���r������[�9lH�+��d���O"���T�E"��T�7'3W��B#n9Pe�x6"��c$���\���F�"Iz�z����84��R��IQ%��Fun���g�4�I'Dے�!M<���
�kz~OO�;w�����'7�xN1 BBޒH1����0�n%�~9_n�b�M� �!EQE<��T��ԱR�-hZQJ(��QJ���R6�pa�Ih�̄�@�I$�a)�!(0�U0%dDуA���A(DP��X௹���|;w%�%�q�a�K�.�]�ƈ!����7�B�c-J�Q����7���=��(�MG�yR���h��5y��xǎ�[���4w)>Rİ�6�°��6����,>g��N�?˓��DO�rd��bX�uY8�)@�s@���q/L�����mci%Ա]�y鯰��9Q���;^�rQcG�ڰ���������Ab�8�iF�cE�,��g����j~ަ����*J�*TJ�m�8�7�z'�pl�`YE�%Ҍ����>����dn`�X�D��Z=��ǥ�w��&o�:c�9�`N�{yݍg7D�?�����4�=x�k9H�sG����	������r7�LjH��=��b�=K<.��ԭfN�Ԛ��#О�81g~��$I,6=+�.y�:c�IsR�P�/p�Acq��@��F�C�#j���%����ˡ%Rܝ(����N���ZR}�{��v�{��O������usVE�qF��դY��F�3\�)��*T��u4D�=Y��&V+��3�Gs���k����Нy�L�^(��J���uys�7&���:�52�͆C��-���5pM�c��Yœz��z��%��qө�C7z��a��>�$a�\))���I���&��Y�V�]6�>Lj�������=,KMQ���"�(H2�&� 