BZh91AY&SY�)� �߀Py���g߰����`	_<��:r C�: �2���(�i�@h    S@"�M��Ѡ4  h4��P        MHI�SA�2 2 @ �101��&"��#B=2�F��ML�FMM�����Ag�	D����Qn����w4�B�� _
�ER�ujf^BI�HFI&!2fi��N�_{x�8j�kUTUUE��j��eQU�      pP` ��reG�"�Dd�0��A��]��t�y�:���'���)x̽��.'�飯z����s!^B��R����j����"*"n����?����нv�c{��5�}{LC��U=Kǵ���!^B�����rY� ��F�h����� f`b����f��d�}V	��79�?<?�[�uw�6�F�����޳jf�Nswwy��33F����ڪ��(�>O{��0�2�����A�|�\;2�=�Hi�S}ĕ��F�,R�	hr^A4�$��u��F�v`�<h��y����-\�EYd��R��p^�c�5Ӈ�`a�)"�Ch�t7 V����1�ɒ��T@�qA�ۚ�f��@�u����8�iR&t�.�Ɠ���� ON��χ~|k�I&E*��HG�׹@B-nq7DB1�j�K(q"j-���LM�8�xG)�Cw�F�$�.��vm a�]MÛWF`�U��Zx$�oB�M��i���k�Q\��s�9��l6Ԟ���;��/)�\�����|I$�V����egOAg�đ�R�!��0�����|�餻�,�GԜ��g�n����v1^,��RI$�|���i�9��9h��0<�(�n@�(���������*��^꠪ͭI$���S����
���q"&��3s��AQ����o^""
I$��i+g��D��p����|5�4�+�A%�o䓛މ���-���4�婦q�^��}��Ii,���6��:#,UڭW����7�X���K�0��Ȉ��ăY�4W\:�
�ASfS�P��G	8{���b�j,Q�>"g�{ʂ��A�^��0�e/�\Rh��	:*I$P�B��LFԔ`�����DA� �0�D� �b���i%KZ�h�J�AVcbŤ��4梤��k�;�@�,�t:0#�d6�>�LkjR�n��<P4��Հ�#c).�i�Ő�|�>����D�w�j;�Je���;=�����6�Q�6=�^�N����;��k9�PC��!�G�8lzH=f���Ty�$��χ؃¡�����x�.�P�;��(���w�=S��-�H�V�����<>�p_���d��^�l��C���G������z@���Ia�6��2\I��'�^(lN~�R\��(L���00$Ne�
�,n	�7v!�~qC6a�`lj0H�&��{\E
?//��87[$��Q��$/[&��*'@*�D���%���
H%!�^,����=IT� ���5}������CY� "��;ͭ���a�np
���IԄ�9�#C��<W& �[��q^t�b�A#'2�J�	m�%�Vm���h�$!�c�MA������P����u��+Q"NߗٽX���z���G[$�:ͅ����lnry:d4���r�0t�G�E��s�wb85U"i$�#t���C�������������������DB�CP�P�P��#��Xu'��q��"�3�SE�h��.�'I9����8Q/���^V�U��<��F�7&ˢ
�2f�q�M����]��y���p"��Yp2����������V"v��)K�r�~�&���:�!
p``���ܑN$��m�