BZh91AY&SY�ק� �_�Py���g߰����`>���>����  ϵ(([pZP�I�'�xQ��    @��hJI�@��20�i�� aO{�U h��M�Mh�  Jz�f�
�i�2i� �    "�m!���4CM  �$���xQ<OT�bO(Ѡ�hjz������D���>ᐙQn���.��|�R�����U��R/~� 8�8u�qꦛ���MH��P	(�Je ��	��UMR3ET�~�wC�����5.���3 7*����Ώ�r����ZnD����ƤS���:�uJ��Y�M/g�3�u
��C\ˈg/�6N�ʫ!j�,�g�o8L�{	�j����X3H�b����ۋhDQ��`�%�Z�h���ՍE�]�x����V4z���G<0AA�h�s��0Wo�p	�=z���|��P�*�����T��U^���IU�Zt�A2���*�If[5�$�H��Ī�0��z<��pq�d�f���zA�,��)T����m��|�*���|F�ǃY��SKqisB�2m�1D�a�֡��8��c�wc��b����gk�-��Ȯe=8�����u�b7��E�Ѳ��.''��N�bRd�\$K���!m<=�7s�-�ؚ�%�w�Y"�nKxjf�LoRkRs�-�Ama;ղ�LZ�:o�՛����Sp�8dè�`����^f3>Q�g�"#�'^��]3�s�u훾�ob��r�L̲�B�� '}�M�Ƕ�8�͸���<�c�M.�9`\ӊ;e�4Ù&����ɶ(��U�ش�3tLE���1���1Q/,�lJ��2TN�Sr��`z89���g�kB�d�G���0��I$�7w�ڊ�Ǒ<�1V��`�`����]��1M��(f�xz��"�Mi��C1�ˀq�P����!Lco�8I$�e��=[A����w��]��`l��)��6k&�h�T��'��ƧV�;�0�^ݦ�a�G��n�_h�Q$�I�"��-��k96�ĕ]q�\�Ikc��L'\='8�&����i�4\[��Z����3��EH1��|��I$�ºH�j�����$�s�c����2���z��m뗀�����Њ��5��^�Ȓ�9�k	�@JKM���.��qX!��I&V)5�]3�#�<�,�g##�hPs�S�*a����^�c˼ᇗ����I�6�T$��*ghN��GN��61K���`HWc#�k"���#(f�z5Hn�n��Qg�\2��%�-���5���[� D4�`�
�6��5S��Y'����V1�
�b��ܷ�37�ݎ~��ԯC��M�:b��:��w�{��,""I��Q��h���u�^�g��Q����b���\r���*� �JH�"@�H��h� E� ���0S"!kQ�j�H��kE�V���KP�q��CQ����:���AI�I�$<+B���~�Ze��_v��v�wР�����qB��NU�,v�.N�`2�:+E�.� 9_yQ�-����7�̃���Q�'��^Û�~Md)0��I	��G���i�C���aa(���H.�d���T~�r��h#hm��Iڞ@�r�;��tIA�D�b�?F�QG����� �('��-Z�x���+n�0�~�RsQ0�C:"A��Ҹ��vPGe�#E�3�v�v�\�#Ȟ=n����Ō@�$�%or�y�$���{�5j:�G{h�Ѱ�1�+�zh#=ޞ��6���*���A�L�'Q�h�����z�fL�/z�>`��/AC����V��pQQikU�](������<�$����Ux*�a܄|󞄱�-k�l��o$�,S���`�se��W Qb�uXq���6�yq�����QS�V �۠��7̏a�D3%(K�hY8�
����تV"U�j�m����X8a~�	���D����"K����1&ǁ�fìw4-a���h9�	��A��Gq�<��ܪ*�*���*�������,**(��������*��������#

"�*�(��
�(�������A
�+�1I��t��@�0I�25k	3��bx�4��b*fE�;
g�@���>#t�UG#�6'!|!D�zc��.��Cs��͇�#35�ĆQ��k.�%C�D�����Aը�F��"p�����/��1��=S�A��G�.�p�!_�Op